library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",X"00",
		X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",X"00",
		X"11",X"99",X"DD",X"DD",X"FF",X"77",X"33",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"33",X"22",X"00",X"44",X"66",X"77",X"55",X"44",X"44",X"00",X"00",
		X"44",X"FF",X"FF",X"44",X"44",X"CC",X"CC",X"00",X"00",X"77",X"77",X"66",X"33",X"11",X"00",X"00",
		X"EE",X"FF",X"11",X"11",X"11",X"33",X"22",X"00",X"00",X"55",X"55",X"55",X"55",X"77",X"77",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"00",X"44",X"44",X"44",X"66",X"33",X"11",X"00",
		X"00",X"00",X"88",X"FF",X"77",X"00",X"00",X"00",X"66",X"77",X"55",X"44",X"44",X"66",X"66",X"00",
		X"66",X"77",X"DD",X"DD",X"99",X"99",X"66",X"00",X"00",X"33",X"44",X"44",X"55",X"77",X"33",X"00",
		X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"FF",X"FF",X"44",X"44",X"44",X"FF",X"FF",X"00",X"11",X"33",X"66",X"44",X"66",X"33",X"11",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"77",X"00",
		X"22",X"33",X"11",X"11",X"33",X"EE",X"CC",X"00",X"22",X"66",X"44",X"44",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"33",X"11",X"11",X"FF",X"FF",X"00",X"11",X"33",X"66",X"44",X"44",X"77",X"77",X"00",
		X"11",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",X"44",X"44",X"44",X"44",X"77",X"77",X"00",X"00",
		X"00",X"88",X"88",X"88",X"88",X"FF",X"FF",X"00",X"44",X"44",X"44",X"44",X"44",X"77",X"77",X"00",
		X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"03",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C8",X"C8",X"CC",X"CC",X"EE",X"AA",X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"33",
		X"9B",X"DD",X"FF",X"F7",X"79",X"F1",X"C0",X"00",X"33",X"30",X"70",X"61",X"10",X"00",X"00",X"00",
		X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"10",X"10",X"11",X"11",X"33",X"33",
		X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"77",X"77",X"DD",X"FF",X"FF",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"EE",X"00",X"DD",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"00",X"EE",X"DD",X"00",X"00",
		X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"33",X"77",X"77",X"33",X"11",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"11",X"33",X"77",X"77",X"33",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"88",
		X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"EE",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"77",
		X"33",X"33",X"33",X"33",X"FF",X"EE",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"FF",X"77",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"00",X"88",X"44",X"22",X"00",X"88",X"44",X"22",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"88",X"22",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"33",X"00",X"00",X"00",
		X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"EE",X"22",X"22",X"00",X"11",X"22",X"22",X"22",X"33",
		X"AA",X"AA",X"AA",X"22",X"00",X"00",X"00",X"EE",X"22",X"22",X"22",X"11",X"00",X"22",X"22",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",
		X"33",X"33",X"77",X"77",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"33",X"33",X"77",X"77",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",X"33",X"33",X"33",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",
		X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"EE",X"EE",X"EE",X"66",X"22",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FF",X"BB",X"BB",X"33",X"33",X"FF",X"EE",X"DD",X"DD",X"DD",X"DD",X"CC",X"CC",X"FF",X"77",
		X"33",X"33",X"BB",X"BB",X"BB",X"FF",X"FF",X"00",X"CC",X"CC",X"DD",X"DD",X"DD",X"FF",X"FF",X"CC",
		X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"77",X"FF",X"CC",X"CC",X"66",X"FF",X"FF",X"CC",
		X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"EE",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"77",
		X"00",X"EE",X"FF",X"33",X"33",X"33",X"FF",X"FF",X"00",X"77",X"FF",X"CC",X"CC",X"CC",X"FF",X"77",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",X"CC",X"CC",X"FF",X"FF",
		X"00",X"88",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"00",X"77",X"FF",X"CC",X"CC",X"CC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"0C",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"CC",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"77",X"88",X"88",X"77",X"00",X"99",X"AA",X"AA",
		X"3E",X"3E",X"DE",X"1E",X"DE",X"3E",X"3E",X"DE",X"C7",X"C7",X"B7",X"87",X"B7",X"C7",X"C7",X"B7",
		X"F0",X"1E",X"1E",X"9E",X"9E",X"1E",X"1E",X"DE",X"F0",X"87",X"87",X"97",X"97",X"87",X"87",X"B7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"20",X"90",X"80",X"00",X"00",X"30",X"30",X"10",X"10",X"00",X"00",
		X"41",X"21",X"12",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"0C",X"8C",X"0C",X"00",X"00",X"00",X"07",X"0F",X"0F",X"C3",X"1F",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"08",X"0F",X"2F",X"4F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"07",X"4F",X"0F",X"A7",X"87",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"D3",X"87",X"97",X"0F",X"2F",X"07",X"00",X"00",X"33",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"08",X"0E",X"8E",X"1F",X"0F",
		X"0C",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"4F",X"1F",X"0F",X"4F",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"01",X"03",X"87",X"87",X"87",X"47",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"10",
		X"EF",X"47",X"07",X"07",X"03",X"01",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"00",
		X"00",X"FF",X"FF",X"08",X"00",X"88",X"CC",X"77",X"00",X"00",X"11",X"33",X"33",X"11",X"13",X"00",
		X"33",X"88",X"00",X"00",X"88",X"FF",X"77",X"00",X"11",X"11",X"33",X"33",X"13",X"11",X"00",X"00",
		X"00",X"00",X"26",X"EE",X"CC",X"00",X"CC",X"CC",X"00",X"8C",X"EE",X"66",X"11",X"77",X"CC",X"00",
		X"CC",X"00",X"88",X"CE",X"66",X"22",X"00",X"00",X"CC",X"7F",X"33",X"00",X"6E",X"CC",X"88",X"00",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"20",
		X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"10",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"0C",X"0F",X"CF",X"2F",X"0F",X"0F",
		X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"44",X"54",X"32",
		X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"30",X"F0",X"F0",X"F0",X"F0",
		X"68",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"F0",X"C3",X"F0",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"0F",X"0F",X"0D",X"02",X"01",X"00",X"00",X"01",X"05",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"08",X"0E",X"0F",X"2F",X"17",
		X"8C",X"0C",X"0C",X"0C",X"0C",X"08",X"00",X"00",X"0B",X"05",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"F1",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"20",
		X"E0",X"F1",X"E0",X"E0",X"00",X"00",X"00",X"00",X"20",X"20",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"DD",
		X"22",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"0F",X"0F",X"FF",X"FF",X"0F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"0F",X"CF",X"FF",X"0F",X"0F",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"CF",X"3F",X"FF",X"FF",X"3F",X"0F",X"0F",X"0F",X"0F",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"C3",X"F0",X"0F",X"0F",X"F0",X"0F",X"0F",X"C3",X"F0",X"F0",
		X"F0",X"F0",X"0F",X"0F",X"C3",X"F0",X"3C",X"0F",X"F0",X"0F",X"0F",X"C3",X"3C",X"0F",X"C3",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"3C",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"00",X"33",X"74",X"74",X"F8",X"F9",X"F9",X"F9",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"FF",X"F9",X"F9",X"F9",X"F8",X"74",X"74",X"33",X"00",
		X"FF",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"FF",
		X"00",X"CC",X"E2",X"E2",X"F1",X"F9",X"F9",X"F9",X"FF",X"F0",X"F0",X"FE",X"11",X"00",X"00",X"00",
		X"F9",X"F9",X"F9",X"F1",X"E2",X"E2",X"CC",X"00",X"00",X"00",X"00",X"11",X"FE",X"F0",X"F0",X"FF",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FF",X"F0",X"F0",X"FE",X"11",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"11",X"FE",X"F0",X"F0",X"FF",
		X"FF",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"FF",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E2",X"E2",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"E2",X"E2",X"CC",X"00",
		X"00",X"33",X"74",X"74",X"F8",X"F8",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"F8",X"F8",X"74",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"33",X"74",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E2",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F8",X"F8",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F9",X"F8",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F1",X"F1",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F9",X"F1",X"F1",X"FF",X"00",X"00",X"00",X"00",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F1",
		X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"11",X"FE",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"FE",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"74",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"E2",X"F1",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"F7",X"F0",X"F0",X"F0",X"F9",X"F9",X"F9",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F0",X"F0",X"F0",X"F7",X"88",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"F8",X"F8",X"F9",X"F9",X"F9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"0C",X"0C",X"8C",X"0C",X"00",X"00",X"30",X"30",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"20",X"90",X"80",X"00",X"00",X"00",X"07",X"0F",X"0F",X"C3",X"1F",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"41",X"21",X"12",X"03",X"03",X"01",X"00",X"00",X"07",X"08",X"0F",X"2F",X"4F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"00",X"07",X"4F",X"0F",X"A7",X"87",X"00",X"00",X"00",X"08",X"0E",X"8E",X"1F",X"0F",
		X"0C",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"33",X"10",X"10",X"10",X"00",X"00",X"00",X"00",
		X"D3",X"87",X"97",X"0F",X"2F",X"07",X"00",X"00",X"4F",X"1F",X"0F",X"4F",X"0E",X"08",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"10",
		X"00",X"00",X"01",X"03",X"87",X"87",X"87",X"47",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"47",X"07",X"07",X"03",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"00",
		X"00",X"00",X"26",X"EE",X"CC",X"00",X"CC",X"CC",X"00",X"00",X"11",X"33",X"33",X"11",X"13",X"00",
		X"00",X"FF",X"FF",X"08",X"00",X"88",X"CC",X"77",X"00",X"8C",X"EE",X"66",X"11",X"77",X"CC",X"00",
		X"CC",X"00",X"88",X"CE",X"66",X"22",X"00",X"00",X"11",X"11",X"33",X"33",X"13",X"11",X"00",X"00",
		X"33",X"88",X"00",X"00",X"88",X"FF",X"77",X"00",X"CC",X"7F",X"33",X"00",X"6E",X"CC",X"88",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"20",
		X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0C",X"0F",X"CF",X"2F",X"0F",X"0F",
		X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"01",X"01",X"00",X"00",X"00",
		X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"44",X"54",X"32",
		X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"00",X"00",X"00",X"30",X"F0",X"F0",X"F0",X"F0",
		X"68",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"C3",X"F0",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"01",X"05",X"02",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"0F",X"0F",X"0D",X"02",X"01",X"00",X"00",X"00",X"08",X"0E",X"0F",X"2F",X"17",
		X"8C",X"0C",X"0C",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"05",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"F8",X"70",X"30",X"10",
		X"00",X"00",X"00",X"0C",X"04",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"07",X"04",X"07",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"02",X"03",X"00",X"00",X"0F",X"00",X"00",X"00",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"04",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"07",X"04",X"07",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",
		X"02",X"03",X"00",X"0D",X"05",X"07",X"00",X"00",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"04",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"07",X"04",X"07",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",
		X"02",X"03",X"00",X"07",X"05",X"0D",X"00",X"00",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"04",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"07",X"04",X"07",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",
		X"02",X"03",X"00",X"0F",X"00",X"00",X"00",X"00",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"03",X"02",X"03",X"00",X"0F",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
		X"01",X"00",X"0F",X"08",X"0F",X"00",X"0C",X"00",X"0F",X"00",X"08",X"08",X"08",X"00",X"00",X"00",
		X"0E",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"03",X"02",X"03",X"00",X"0F",X"01",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"05",X"05",X"00",
		X"0F",X"08",X"0F",X"00",X"04",X"04",X"0C",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"02",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"03",X"02",X"03",X"00",X"0F",X"01",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"05",X"07",X"00",
		X"0F",X"08",X"0F",X"00",X"0C",X"04",X"04",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"0F",
		X"0E",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"55",X"DD",X"DD",X"55",X"55",X"33",
		X"66",X"66",X"55",X"DD",X"DD",X"77",X"77",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"DD",X"DD",X"55",X"55",X"33",
		X"00",X"00",X"00",X"00",X"88",X"88",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"55",X"DD",X"DD",X"55",X"55",X"33",X"00",X"00",X"00",X"00",X"88",X"88",X"44",X"44",
		X"11",X"11",X"55",X"55",X"DD",X"99",X"11",X"DD",X"99",X"CC",X"EE",X"BB",X"99",X"CC",X"EE",X"BB",
		X"AA",X"88",X"AA",X"AA",X"BB",X"99",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",
		X"11",X"11",X"11",X"DD",X"11",X"FF",X"00",X"00",X"99",X"CC",X"EE",X"BB",X"99",X"FF",X"CC",X"88",
		X"99",X"BB",X"99",X"88",X"88",X"FF",X"00",X"00",X"EE",X"22",X"EE",X"77",X"00",X"FF",X"00",X"00",
		X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"CC",X"EE",X"BB",X"99",X"CC",X"EE",X"BB",
		X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"DD",X"11",X"99",X"CC",X"EE",X"BB",X"99",X"CC",X"EE",X"BB",
		X"88",X"88",X"88",X"88",X"AA",X"AA",X"BB",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"88",X"88",X"88",X"CC",X"44",X"44",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"DD",X"DD",X"DD",X"55",X"55",X"77",X"33",
		X"66",X"66",X"55",X"55",X"DD",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"11",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"33",X"FF",X"55",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"77",X"33",X"33",X"33",X"11",X"11",X"CC",X"44",X"44",X"66",X"66",X"66",X"77",X"55",
		X"CC",X"99",X"BB",X"EE",X"CC",X"99",X"BB",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"99",X"BB",X"EE",X"DD",X"BB",X"BB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"99",X"BB",X"EE",X"CC",X"99",X"BB",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"99",X"BB",X"EE",X"CC",X"99",X"BB",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",X"FF",X"FF",X"77",X"77",
		X"00",X"11",X"11",X"11",X"33",X"FF",X"FF",X"FF",X"88",X"88",X"88",X"88",X"88",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"33",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"77",X"00",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"77",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"00",X"CC",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"33",X"33",X"77",X"77",X"77",
		X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"EE",X"EE",X"EE",X"FF",X"FF",X"FF",X"77",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"00",X"E0",X"C0",X"80",X"C0",X"E0",X"E0",X"80",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",
		X"00",X"10",X"F0",X"F0",X"F0",X"F3",X"F3",X"F0",X"00",X"F0",X"F1",X"F2",X"F2",X"F1",X"F1",X"F2",
		X"80",X"E0",X"E0",X"C0",X"80",X"C0",X"E0",X"00",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"00",
		X"F0",X"F3",X"F3",X"F0",X"F0",X"F0",X"10",X"00",X"F2",X"F1",X"F1",X"F2",X"F2",X"F1",X"F0",X"00",
		X"00",X"C0",X"E0",X"E0",X"C0",X"80",X"C0",X"E0",X"00",X"00",X"00",X"10",X"30",X"30",X"70",X"70",
		X"00",X"10",X"F0",X"F0",X"F0",X"F3",X"F3",X"F0",X"00",X"F0",X"F1",X"F2",X"F2",X"F1",X"F1",X"F2",
		X"E0",X"C0",X"80",X"C0",X"E0",X"E0",X"C0",X"00",X"70",X"70",X"30",X"30",X"10",X"00",X"00",X"00",
		X"F0",X"F3",X"F3",X"F0",X"F0",X"F0",X"10",X"00",X"F2",X"F1",X"F1",X"F2",X"F2",X"F1",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"11",X"33",X"77",X"77",X"33",X"11",
		X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"77",X"33",X"11",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"BC",X"3C",X"0F",X"8F",X"FF",X"FF",X"00",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"BC",X"3C",X"0F",X"8F",X"FF",X"FF",X"11",X"00",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"BC",X"3C",X"0F",X"8F",X"FF",X"FF",X"00",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"BC",X"3C",X"0F",X"8F",X"FF",X"FF",X"11",X"00",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"CF",X"8F",X"8F",X"CF",X"FF",X"00",X"FF",X"FF",X"7F",X"F3",X"F3",X"7F",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"CF",X"8F",X"8F",X"CF",X"FF",X"11",X"00",X"FF",X"7F",X"F3",X"F3",X"7F",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"CF",X"8F",X"8F",X"CF",X"FF",X"00",X"FF",X"FF",X"7F",X"F3",X"F3",X"7F",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"CF",X"8F",X"8F",X"CF",X"FF",X"11",X"00",X"FF",X"7F",X"F3",X"F3",X"7F",X"FF",X"FF",X"00",
		X"00",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"11",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"11",X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"77",X"33",X"33",X"11",X"00",X"00",X"00",
		X"FF",X"FF",X"8F",X"0F",X"3C",X"BC",X"11",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"00",
		X"00",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"88",X"00",X"00",X"00",X"01",X"30",X"30",X"67",X"77",
		X"00",X"11",X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"77",X"67",X"30",X"30",X"01",X"00",X"00",X"00",
		X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"CC",X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"00",X"00",X"00",X"01",X"30",X"30",X"67",X"77",
		X"00",X"11",X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"CC",X"00",X"77",X"67",X"30",X"30",X"01",X"00",X"00",X"00",
		X"FF",X"3F",X"1F",X"1F",X"3F",X"FF",X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"06",X"02",X"0C",X"00",X"02",X"02",X"0A",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"0F",X"04",X"02",X"01",X"02",X"0C",X"00",X"08",X"0E",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"02",X"0C",X"00",X"0C",X"02",X"02",X"02",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"09",X"09",X"09",X"07",X"00",X"0F",X"0C",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"11",X"33",X"33",X"77",X"77",X"88",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"77",X"77",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"88",X"88",
		X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"33",
		X"10",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"C0",X"E6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"33",X"30",X"70",X"61",X"10",X"00",X"00",X"00",
		X"DD",X"DD",X"DD",X"F7",X"79",X"F1",X"C0",X"00",X"FF",X"FF",X"DD",X"FF",X"FF",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"EE",X"00",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"20",X"62",X"EE",X"EE",X"00",X"00",X"00",X"00",X"20",X"32",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"33",X"30",X"70",X"61",X"10",X"00",X"00",X"00",
		X"22",X"9B",X"DD",X"F7",X"79",X"F1",X"C0",X"00",X"33",X"77",X"DD",X"FF",X"FF",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"33",X"FF",X"FB",X"FF",X"77",X"77",X"33",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"FE",X"00",X"00",X"00",X"10",X"61",X"70",X"30",X"33",
		X"00",X"C0",X"F1",X"79",X"F7",X"FF",X"88",X"FF",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"77",X"FF",
		X"FC",X"FE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"00",X"00",X"00",
		X"FF",X"FF",X"BB",X"FF",X"FF",X"FF",X"33",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",
		X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"61",X"70",X"30",X"33",
		X"00",X"C0",X"F1",X"79",X"E6",X"CC",X"9B",X"EE",X"00",X"00",X"FE",X"EC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"00",X"00",X"00",
		X"CC",X"EE",X"BB",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"00",X"88",X"CC",X"EC",X"FE",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"10",X"61",X"70",X"30",X"33",
		X"00",X"C0",X"F1",X"79",X"F7",X"EE",X"CD",X"FF",X"00",X"00",X"EE",X"FF",X"FF",X"77",X"CC",X"00",
		X"00",X"00",X"00",X"C0",X"CC",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"00",X"00",X"00",
		X"CC",X"FF",X"BB",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"EE",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"00",X"00",X"00",X"10",X"61",X"70",X"30",X"33",
		X"00",X"C0",X"F1",X"79",X"F7",X"FF",X"DD",X"9B",X"00",X"00",X"EE",X"FF",X"FF",X"DD",X"77",X"77",
		X"EE",X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"00",X"00",X"00",
		X"AA",X"EE",X"CC",X"CC",X"C8",X"C8",X"00",X"00",X"33",X"33",X"11",X"11",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"11",X"33",X"30",X"00",X"00",X"00",
		X"00",X"77",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"DD",X"FF",X"33",
		X"CC",X"C0",X"E0",X"68",X"80",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"11",X"00",X"00",X"00",
		X"00",X"33",X"EE",X"FF",X"FF",X"77",X"00",X"00",X"FF",X"3B",X"77",X"FE",X"E9",X"F8",X"30",X"00",
		X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"33",
		X"00",X"00",X"C8",X"C8",X"CC",X"CC",X"EE",X"AA",X"00",X"00",X"10",X"10",X"11",X"11",X"33",X"33",
		X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"33",X"30",X"70",X"61",X"10",X"00",X"00",X"00",
		X"9B",X"DD",X"FF",X"F7",X"79",X"F1",X"C0",X"00",X"77",X"77",X"DD",X"FF",X"FF",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"10",X"61",X"70",X"30",X"33",
		X"00",X"C0",X"F1",X"79",X"F7",X"EE",X"CD",X"FF",X"00",X"00",X"EE",X"FF",X"FF",X"77",X"CC",X"00",
		X"00",X"00",X"00",X"C0",X"CC",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"00",X"00",X"00",
		X"CC",X"FF",X"BB",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"EE",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"00",X"00",X"00",X"10",X"61",X"70",X"30",X"33",
		X"00",X"C0",X"F1",X"79",X"F7",X"FF",X"DD",X"9B",X"00",X"00",X"EE",X"FF",X"FF",X"DD",X"77",X"77",
		X"EE",X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"00",X"00",X"00",
		X"AA",X"EE",X"CC",X"CC",X"C8",X"C8",X"00",X"00",X"33",X"33",X"11",X"11",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"11",X"33",X"30",X"00",X"00",X"00",
		X"00",X"77",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"DD",X"FF",X"33",
		X"CC",X"C0",X"E0",X"68",X"80",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"11",X"00",X"00",X"00",
		X"00",X"33",X"EE",X"FF",X"FF",X"77",X"00",X"00",X"FF",X"3B",X"77",X"FE",X"E9",X"F8",X"30",X"00",
		X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"11",X"11",X"33",X"33",X"33",
		X"00",X"00",X"C8",X"C8",X"CC",X"CC",X"EE",X"AA",X"00",X"00",X"10",X"10",X"11",X"11",X"33",X"33",
		X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"00",X"33",X"30",X"70",X"61",X"10",X"00",X"00",X"00",
		X"9B",X"DD",X"FF",X"F7",X"79",X"F1",X"C0",X"00",X"77",X"77",X"DD",X"FF",X"FF",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"10",X"61",X"70",X"30",X"33",
		X"00",X"C0",X"F1",X"79",X"F7",X"EE",X"CD",X"FF",X"00",X"00",X"EE",X"FF",X"FF",X"77",X"CC",X"00",
		X"00",X"00",X"00",X"C0",X"CC",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"00",X"00",X"00",
		X"CC",X"FF",X"BB",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"EE",X"00",
		X"00",X"00",X"00",X"88",X"CC",X"CC",X"EE",X"EE",X"00",X"00",X"00",X"10",X"61",X"70",X"30",X"33",
		X"00",X"C0",X"F1",X"79",X"F7",X"FF",X"DD",X"9B",X"00",X"00",X"EE",X"FF",X"FF",X"DD",X"77",X"77",
		X"EE",X"EE",X"EE",X"CC",X"CC",X"88",X"00",X"00",X"33",X"33",X"33",X"11",X"11",X"00",X"00",X"00",
		X"AA",X"EE",X"CC",X"CC",X"C8",X"C8",X"00",X"00",X"33",X"33",X"11",X"11",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"11",X"33",X"30",X"00",X"00",X"00",
		X"00",X"77",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"DD",X"FF",X"33",
		X"CC",X"C0",X"E0",X"68",X"80",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"11",X"00",X"00",X"00",
		X"00",X"33",X"EE",X"FF",X"FF",X"77",X"00",X"00",X"FF",X"3B",X"77",X"FE",X"E9",X"F8",X"30",X"00",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"CC",X"00",X"00",X"11",X"33",X"30",X"00",X"00",X"00",
		X"00",X"77",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"DD",X"FF",X"33",
		X"CC",X"C0",X"E0",X"68",X"80",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"11",X"00",X"00",X"00",
		X"00",X"33",X"EE",X"FF",X"FF",X"77",X"00",X"00",X"FF",X"3B",X"77",X"FE",X"E9",X"F8",X"30",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
