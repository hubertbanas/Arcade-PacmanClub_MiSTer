library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"3E",X"00",X"C3",X"D5",X"1F",X"00",X"00",X"77",X"23",X"10",X"FC",X"C9",X"C3",X"65",X"09",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"78",X"87",X"D7",X"5F",X"23",X"56",X"EB",X"C9",
		X"E1",X"87",X"D7",X"5F",X"23",X"56",X"EB",X"E9",X"E1",X"46",X"23",X"4E",X"23",X"E5",X"18",X"12",
		X"11",X"90",X"4C",X"06",X"10",X"C3",X"51",X"00",X"C3",X"19",X"2F",X"50",X"32",X"07",X"50",X"C3",
		X"38",X"00",X"2A",X"80",X"4C",X"70",X"2C",X"71",X"2C",X"20",X"02",X"2E",X"C0",X"22",X"80",X"4C",
		X"C9",X"1A",X"A7",X"28",X"06",X"1C",X"1C",X"1C",X"10",X"F7",X"C9",X"E1",X"06",X"03",X"7E",X"12",
		X"23",X"1C",X"10",X"FA",X"E9",X"00",X"C3",X"D9",X"B6",X"C3",X"FA",X"1E",X"32",X"C0",X"50",X"31",
		X"C0",X"4F",X"AF",X"21",X"00",X"50",X"01",X"08",X"08",X"CF",X"21",X"00",X"4C",X"06",X"BE",X"CF",
		X"CF",X"CF",X"CF",X"21",X"40",X"50",X"06",X"40",X"CF",X"32",X"C0",X"50",X"CD",X"68",X"20",X"32",
		X"C0",X"50",X"06",X"00",X"CD",X"46",X"20",X"32",X"C0",X"50",X"21",X"C0",X"4C",X"22",X"80",X"4C",
		X"22",X"82",X"4C",X"3E",X"FF",X"06",X"40",X"CF",X"3E",X"01",X"32",X"00",X"50",X"21",X"74",X"36",
		X"11",X"E8",X"4D",X"01",X"10",X"00",X"ED",X"B0",X"FB",X"2A",X"82",X"4C",X"7E",X"A7",X"FA",X"B9",
		X"00",X"36",X"FF",X"2C",X"46",X"36",X"FF",X"2C",X"20",X"02",X"2E",X"C0",X"22",X"82",X"4C",X"21",
		X"B9",X"00",X"E5",X"E7",X"46",X"20",X"C3",X"22",X"74",X"20",X"62",X"22",X"29",X"23",X"75",X"24",
		X"68",X"20",X"82",X"24",X"52",X"25",X"8E",X"25",X"CB",X"25",X"13",X"26",X"5D",X"26",X"8C",X"26",
		X"BB",X"26",X"EA",X"26",X"0D",X"00",X"8C",X"24",X"B5",X"22",X"6B",X"28",X"D2",X"24",X"8A",X"22",
		X"41",X"20",X"19",X"27",X"1D",X"29",X"90",X"28",X"E4",X"29",X"64",X"2A",X"15",X"96",X"1B",X"2A",
		X"5F",X"24",X"9C",X"24",X"DA",X"2A",X"96",X"28",X"35",X"01",X"C3",X"13",X"24",X"60",X"3E",X"19",
		X"21",X"79",X"37",X"01",X"00",X"71",X"EF",X"AD",X"00",X"71",X"BA",X"24",X"20",X"30",X"C3",X"00",
		X"00",X"C9",X"78",X"21",X"D1",X"31",X"EF",X"AD",X"C9",X"7B",X"BA",X"24",X"38",X"AE",X"66",X"01",
		X"7B",X"01",X"4D",X"83",X"78",X"65",X"56",X"76",X"11",X"60",X"45",X"63",X"67",X"65",X"89",X"76",
		X"78",X"65",X"90",X"78",X"0A",X"79",X"0A",X"79",X"80",X"79",X"89",X"76",X"90",X"78",X"43",X"65",
		X"45",X"7F",X"89",X"6A",X"9A",X"67",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",
		X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"01",X"03",X"04",X"06",X"07",
		X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"14",X"14",X"14",X"14",X"14",X"14",
		X"00",X"00",X"00",X"01",X"03",X"04",X"06",X"08",X"0A",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"12",
		X"13",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"00",X"00",X"00",X"E3",X"DD",X"E5",X"FD",X"E5",
		X"C5",X"47",X"CD",X"CD",X"01",X"7E",X"23",X"A7",X"28",X"0C",X"FD",X"77",X"00",X"DD",X"70",X"00",
		X"FD",X"19",X"DD",X"19",X"18",X"EF",X"C1",X"FD",X"E1",X"DD",X"E1",X"E3",X"C9",X"C5",X"FD",X"21",
		X"00",X"40",X"DD",X"21",X"00",X"44",X"42",X"4B",X"11",X"20",X"00",X"78",X"A7",X"28",X"06",X"FD",
		X"19",X"DD",X"19",X"10",X"FA",X"59",X"FD",X"19",X"DD",X"19",X"11",X"E0",X"FF",X"C1",X"C9",X"CD",
		X"62",X"3A",X"3E",X"0F",X"11",X"1A",X"1B",X"CD",X"AB",X"01",X"49",X"4E",X"44",X"55",X"53",X"54",
		X"52",X"49",X"41",X"40",X"41",X"52",X"47",X"45",X"4E",X"54",X"49",X"4E",X"41",X"00",X"06",X"10",
		X"CD",X"79",X"32",X"3E",X"0F",X"11",X"1C",X"1B",X"CD",X"AB",X"01",X"5C",X"40",X"49",X"4E",X"47",
		X"40",X"4F",X"4A",X"45",X"44",X"41",X"40",X"31",X"39",X"39",X"30",X"00",X"06",X"10",X"CD",X"79",
		X"32",X"3E",X"0F",X"11",X"1E",X"1B",X"CD",X"AB",X"01",X"4E",X"55",X"4D",X"45",X"52",X"4F",X"40",
		X"53",X"45",X"52",X"49",X"45",X"40",X"50",X"41",X"43",X"30",X"30",X"30",X"30",X"00",X"06",X"10",
		X"CD",X"79",X"32",X"21",X"00",X"40",X"06",X"04",X"C9",X"7B",X"03",X"4E",X"4F",X"52",X"4D",X"41",
		X"4C",X"40",X"40",X"40",X"40",X"52",X"41",X"50",X"49",X"44",X"4F",X"40",X"40",X"40",X"40",X"54",
		X"55",X"52",X"42",X"4F",X"2F",X"89",X"2F",X"80",X"78",X"03",X"40",X"40",X"40",X"40",X"40",X"40",
		X"44",X"4F",X"42",X"4C",X"45",X"40",X"43",X"4F",X"4D",X"41",X"4E",X"44",X"4F",X"40",X"40",X"40",
		X"40",X"40",X"40",X"2F",X"89",X"2F",X"80",X"78",X"03",X"40",X"40",X"40",X"40",X"40",X"40",X"44",
		X"4F",X"42",X"4C",X"45",X"40",X"43",X"4F",X"4D",X"41",X"4E",X"44",X"4F",X"40",X"40",X"40",X"40",
		X"40",X"40",X"2F",X"81",X"2F",X"80",X"7B",X"03",X"4E",X"4F",X"52",X"4D",X"41",X"4C",X"40",X"2F",
		X"81",X"2F",X"80",X"3B",X"02",X"52",X"41",X"50",X"49",X"44",X"4F",X"40",X"2F",X"81",X"2F",X"80",
		X"FB",X"00",X"54",X"55",X"52",X"42",X"4F",X"2F",X"81",X"2F",X"80",X"92",X"02",X"54",X"55",X"52",
		X"42",X"4F",X"2F",X"81",X"2F",X"80",X"69",X"03",X"40",X"40",X"40",X"40",X"49",X"4E",X"43",X"45",
		X"52",X"54",X"40",X"59",X"4F",X"55",X"52",X"40",X"4E",X"41",X"4D",X"45",X"40",X"40",X"40",X"2F",
		X"89",X"2F",X"80",X"65",X"03",X"40",X"40",X"53",X"45",X"4C",X"45",X"43",X"54",X"40",X"53",X"50",
		X"45",X"45",X"44",X"40",X"50",X"41",X"43",X"4B",X"4D",X"41",X"4E",X"2F",X"89",X"2F",X"80",X"7D",
		X"03",X"40",X"40",X"40",X"50",X"4F",X"52",X"40",X"46",X"41",X"56",X"4F",X"52",X"40",X"4D",X"41",
		X"53",X"40",X"46",X"49",X"43",X"48",X"41",X"53",X"40",X"2F",X"85",X"2F",X"80",X"7D",X"03",X"40",
		X"40",X"50",X"4F",X"52",X"40",X"46",X"41",X"56",X"4F",X"52",X"40",X"53",X"45",X"4C",X"45",X"43",
		X"43",X"49",X"4F",X"4E",X"45",X"40",X"40",X"2F",X"85",X"2F",X"80",X"92",X"02",X"45",X"58",X"54",
		X"52",X"41",X"40",X"4C",X"49",X"46",X"45",X"2F",X"89",X"2F",X"80",X"92",X"02",X"42",X"4F",X"4E",
		X"55",X"53",X"40",X"4E",X"4F",X"4E",X"45",X"2F",X"81",X"2F",X"80",X"92",X"02",X"32",X"30",X"30",
		X"40",X"40",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"85",X"2F",X"80",X"92",X"02",X"33",X"30",X"30",
		X"40",X"40",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"85",X"2F",X"80",X"92",X"02",X"34",X"30",X"30",
		X"40",X"40",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"85",X"2F",X"80",X"92",X"02",X"35",X"30",X"30",
		X"40",X"40",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"85",X"2F",X"80",X"92",X"02",X"36",X"30",X"30",
		X"40",X"40",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"85",X"2F",X"80",X"92",X"02",X"37",X"30",X"30",
		X"40",X"40",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"85",X"2F",X"80",X"92",X"02",X"38",X"30",X"30",
		X"40",X"40",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"85",X"2F",X"80",X"92",X"02",X"35",X"30",X"30",
		X"30",X"40",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"85",X"2F",X"80",X"10",X"11",X"12",X"13",X"14",
		X"01",X"03",X"04",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"14",
		X"21",X"84",X"4C",X"34",X"23",X"35",X"23",X"11",X"4D",X"04",X"01",X"01",X"04",X"34",X"7E",X"E6",
		X"0F",X"EB",X"BE",X"20",X"13",X"0C",X"1A",X"C6",X"10",X"E6",X"F0",X"12",X"23",X"BE",X"20",X"08",
		X"0C",X"EB",X"36",X"00",X"23",X"13",X"10",X"E5",X"21",X"8A",X"4C",X"71",X"2C",X"7E",X"87",X"87",
		X"86",X"3C",X"77",X"2C",X"7E",X"87",X"86",X"87",X"87",X"86",X"3C",X"77",X"C9",X"06",X"A0",X"0A",
		X"60",X"0A",X"60",X"0A",X"A0",X"21",X"6A",X"4C",X"5E",X"23",X"56",X"D5",X"E1",X"77",X"21",X"90",
		X"4C",X"3A",X"8A",X"4C",X"4F",X"06",X"10",X"7E",X"A7",X"28",X"43",X"E6",X"C0",X"07",X"07",X"B9",
		X"30",X"3C",X"35",X"7E",X"E6",X"3F",X"20",X"36",X"77",X"C5",X"E5",X"2C",X"7E",X"2C",X"46",X"21",
		X"AC",X"04",X"E5",X"E7",X"F1",X"0A",X"D0",X"08",X"8F",X"06",X"87",X"14",X"AF",X"11",X"B4",X"11",
		X"B4",X"04",X"B7",X"04",X"B7",X"04",X"B7",X"04",X"B7",X"04",X"DC",X"B5",X"00",X"67",X"89",X"7F",
		X"47",X"65",X"89",X"67",X"00",X"70",X"B5",X"7A",X"9A",X"78",X"AF",X"79",X"E1",X"C1",X"2C",X"2C",
		X"2C",X"10",X"B4",X"C9",X"EF",X"1C",X"86",X"C9",X"3A",X"6E",X"4E",X"FE",X"99",X"17",X"32",X"06",
		X"50",X"1F",X"D0",X"3A",X"00",X"50",X"47",X"CB",X"00",X"3A",X"66",X"4E",X"17",X"E6",X"0F",X"32",
		X"66",X"4E",X"D6",X"0C",X"CC",X"30",X"05",X"CB",X"00",X"3A",X"67",X"4E",X"17",X"E6",X"0F",X"32",
		X"67",X"4E",X"D6",X"0C",X"C2",X"EB",X"04",X"21",X"69",X"4E",X"34",X"CB",X"00",X"3A",X"68",X"4E",
		X"17",X"E6",X"0F",X"32",X"68",X"4E",X"D6",X"0C",X"C0",X"21",X"69",X"4E",X"34",X"C9",X"3A",X"69",
		X"4E",X"A7",X"C8",X"47",X"3A",X"6A",X"4E",X"5F",X"FE",X"00",X"C2",X"15",X"05",X"3E",X"01",X"32",
		X"07",X"50",X"CD",X"30",X"05",X"7B",X"FE",X"08",X"C2",X"1F",X"05",X"AF",X"32",X"07",X"50",X"1C",
		X"7B",X"32",X"6A",X"4E",X"D6",X"10",X"C0",X"32",X"6A",X"4E",X"05",X"78",X"32",X"69",X"4E",X"C9",
		X"3A",X"6B",X"4E",X"21",X"6C",X"4E",X"34",X"96",X"C0",X"77",X"3A",X"6D",X"4E",X"21",X"6E",X"4E",
		X"86",X"27",X"D2",X"47",X"05",X"3E",X"99",X"FE",X"02",X"38",X"12",X"F5",X"C5",X"D5",X"E5",X"3A",
		X"03",X"4E",X"FE",X"01",X"20",X"03",X"EF",X"20",X"0B",X"E1",X"D1",X"C1",X"F1",X"77",X"21",X"9C",
		X"4E",X"CB",X"CE",X"C9",X"21",X"CE",X"4D",X"34",X"7E",X"E6",X"0F",X"20",X"1F",X"7E",X"0F",X"0F",
		X"0F",X"0F",X"47",X"3A",X"D6",X"4D",X"2F",X"B0",X"4F",X"3A",X"6E",X"4E",X"D6",X"01",X"30",X"02",
		X"AF",X"4F",X"28",X"01",X"79",X"AF",X"32",X"05",X"50",X"32",X"04",X"50",X"DD",X"21",X"D8",X"43",
		X"FD",X"21",X"C5",X"43",X"3A",X"00",X"4E",X"FE",X"03",X"CA",X"AB",X"05",X"3A",X"03",X"4E",X"FE",
		X"02",X"D2",X"AB",X"05",X"CD",X"D0",X"05",X"CD",X"DD",X"05",X"C9",X"3A",X"09",X"4E",X"A7",X"3A",
		X"CE",X"4D",X"C2",X"C0",X"05",X"CB",X"67",X"CC",X"D0",X"05",X"C4",X"EA",X"05",X"C3",X"C8",X"05",
		X"CB",X"67",X"CC",X"DD",X"05",X"C4",X"F7",X"05",X"3A",X"70",X"4E",X"A7",X"CC",X"F7",X"05",X"C9",
		X"DD",X"36",X"00",X"50",X"DD",X"36",X"01",X"55",X"DD",X"36",X"02",X"31",X"C9",X"FD",X"36",X"00",
		X"50",X"FD",X"36",X"01",X"55",X"FD",X"36",X"02",X"32",X"C9",X"DD",X"36",X"00",X"40",X"DD",X"36",
		X"01",X"40",X"DD",X"36",X"02",X"40",X"C9",X"FD",X"36",X"00",X"40",X"FD",X"36",X"01",X"40",X"FD",
		X"36",X"02",X"40",X"C9",X"C9",X"3A",X"06",X"4E",X"D6",X"05",X"D8",X"2A",X"08",X"4D",X"06",X"08",
		X"0E",X"10",X"7D",X"32",X"06",X"4D",X"32",X"D2",X"4D",X"91",X"32",X"02",X"4D",X"32",X"04",X"4D",
		X"7C",X"80",X"32",X"03",X"4D",X"32",X"07",X"4D",X"91",X"32",X"05",X"4D",X"32",X"D3",X"4D",X"C9",
		X"3A",X"00",X"4E",X"E6",X"03",X"E7",X"3E",X"06",X"6A",X"06",X"94",X"06",X"EF",X"08",X"3A",X"01",
		X"4E",X"E6",X"01",X"E7",X"48",X"06",X"0C",X"00",X"EF",X"00",X"00",X"EF",X"06",X"00",X"EF",X"01",
		X"00",X"EF",X"14",X"00",X"EF",X"18",X"00",X"EF",X"04",X"00",X"EF",X"1E",X"00",X"EF",X"07",X"00",
		X"21",X"01",X"4E",X"34",X"21",X"01",X"50",X"36",X"01",X"C9",X"CD",X"1B",X"2A",X"3A",X"6E",X"4E",
		X"A7",X"28",X"0C",X"AF",X"32",X"04",X"4E",X"32",X"02",X"4E",X"21",X"00",X"4E",X"34",X"C9",X"C3",
		X"9B",X"3D",X"CD",X"EF",X"08",X"C9",X"06",X"1C",X"CD",X"42",X"00",X"F7",X"4A",X"02",X"00",X"21",
		X"02",X"4E",X"34",X"C9",X"3A",X"03",X"4E",X"E6",X"07",X"E7",X"96",X"07",X"AC",X"06",X"8B",X"08",
		X"0C",X"00",X"D5",X"08",X"A6",X"3F",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"AF",X"32",X"FE",X"4D",
		X"32",X"FF",X"4D",X"CD",X"D3",X"07",X"3A",X"70",X"4C",X"E6",X"03",X"E7",X"C4",X"06",X"F4",X"06",
		X"23",X"07",X"5A",X"07",X"3A",X"71",X"4C",X"A7",X"28",X"0B",X"EF",X"20",X"01",X"AF",X"32",X"71",
		X"4C",X"3C",X"32",X"77",X"4C",X"3A",X"00",X"50",X"CB",X"47",X"CA",X"7E",X"07",X"CB",X"57",X"CA",
		X"E8",X"06",X"CB",X"5F",X"CA",X"17",X"07",X"C0",X"32",X"71",X"4C",X"EF",X"20",X"00",X"3E",X"02",
		X"32",X"70",X"4C",X"C9",X"3A",X"71",X"4C",X"A7",X"28",X"0B",X"EF",X"20",X"02",X"AF",X"32",X"71",
		X"4C",X"3C",X"32",X"77",X"4C",X"3A",X"00",X"50",X"CB",X"47",X"CA",X"7E",X"07",X"CB",X"4F",X"28",
		X"3E",X"CB",X"57",X"CA",X"E8",X"06",X"C0",X"32",X"71",X"4C",X"EF",X"20",X"00",X"3E",X"01",X"32",
		X"70",X"4C",X"C9",X"3A",X"71",X"4C",X"A7",X"28",X"15",X"EF",X"20",X"03",X"3A",X"6E",X"4E",X"FE",
		X"02",X"38",X"03",X"EF",X"20",X"0B",X"AF",X"32",X"71",X"4C",X"3C",X"32",X"77",X"4C",X"3A",X"00",
		X"50",X"CB",X"4F",X"28",X"0A",X"CB",X"47",X"CA",X"7E",X"07",X"CB",X"5F",X"28",X"C9",X"C0",X"32",
		X"71",X"4C",X"EF",X"20",X"00",X"AF",X"32",X"70",X"4C",X"C9",X"3A",X"71",X"4C",X"A7",X"28",X"0B",
		X"EF",X"20",X"0C",X"AF",X"32",X"71",X"4C",X"3C",X"32",X"77",X"4C",X"3A",X"00",X"50",X"CB",X"4F",
		X"CA",X"4F",X"07",X"CB",X"57",X"CA",X"E8",X"06",X"CB",X"5F",X"CA",X"17",X"07",X"C0",X"08",X"3A",
		X"6E",X"4E",X"FE",X"02",X"D8",X"08",X"32",X"71",X"4C",X"EF",X"20",X"00",X"EF",X"20",X"0B",X"3E",
		X"03",X"32",X"70",X"4C",X"C9",X"C9",X"3E",X"00",X"32",X"70",X"4C",X"32",X"71",X"4C",X"32",X"77",
		X"4C",X"AF",X"32",X"72",X"4C",X"CD",X"1B",X"2A",X"EF",X"00",X"01",X"EF",X"01",X"00",X"EF",X"1C",
		X"07",X"EF",X"1C",X"0B",X"EF",X"1E",X"00",X"EF",X"20",X"00",X"EF",X"20",X"07",X"21",X"03",X"4E",
		X"34",X"3E",X"01",X"32",X"D6",X"4D",X"3A",X"71",X"4E",X"FE",X"FF",X"C8",X"EF",X"1C",X"0A",X"EF",
		X"1F",X"00",X"C9",X"CD",X"1B",X"2A",X"3A",X"6E",X"4E",X"FE",X"01",X"06",X"09",X"20",X"0A",X"06",
		X"08",X"18",X"18",X"06",X"37",X"CD",X"DF",X"2A",X"C9",X"FE",X"04",X"D4",X"E3",X"07",X"3A",X"71",
		X"4C",X"A7",X"28",X"05",X"06",X"0B",X"CD",X"DA",X"2A",X"06",X"09",X"CD",X"DF",X"2A",X"3A",X"6E",
		X"4E",X"FE",X"01",X"3A",X"40",X"50",X"28",X"0C",X"CB",X"77",X"20",X"08",X"3E",X"01",X"32",X"70",
		X"4E",X"C3",X"1B",X"08",X"CB",X"6F",X"C0",X"AF",X"32",X"70",X"4E",X"3A",X"6B",X"4E",X"A7",X"28",
		X"48",X"3A",X"77",X"4C",X"A7",X"CA",X"79",X"08",X"3A",X"70",X"4E",X"A7",X"3A",X"6E",X"4E",X"28",
		X"19",X"08",X"3A",X"70",X"4C",X"FE",X"03",X"20",X"0D",X"3A",X"6E",X"4E",X"FE",X"04",X"DA",X"82",
		X"08",X"08",X"C6",X"99",X"27",X"08",X"08",X"C6",X"99",X"27",X"08",X"3A",X"70",X"4C",X"FE",X"03",
		X"20",X"0D",X"3A",X"6E",X"4E",X"FE",X"02",X"DA",X"82",X"08",X"08",X"C6",X"99",X"27",X"08",X"08",
		X"C6",X"99",X"27",X"32",X"6E",X"4E",X"CD",X"1B",X"2A",X"21",X"03",X"4E",X"34",X"AF",X"32",X"D6",
		X"4D",X"3C",X"32",X"CC",X"4E",X"32",X"DC",X"4E",X"C9",X"3E",X"10",X"32",X"BC",X"4E",X"EF",X"20",
		X"0E",X"C9",X"3E",X"04",X"32",X"BC",X"4E",X"EF",X"20",X"0D",X"C9",X"EF",X"00",X"01",X"EF",X"01",
		X"01",X"EF",X"02",X"00",X"EF",X"1C",X"15",X"EF",X"12",X"00",X"EF",X"03",X"00",X"EF",X"1C",X"03",
		X"EF",X"1C",X"06",X"EF",X"29",X"35",X"EF",X"34",X"35",X"EF",X"18",X"00",X"EF",X"1B",X"00",X"AF",
		X"32",X"13",X"4E",X"3A",X"6F",X"4E",X"08",X"3A",X"70",X"4C",X"FE",X"03",X"20",X"04",X"08",X"CB",
		X"27",X"08",X"08",X"32",X"14",X"4E",X"32",X"15",X"4E",X"EF",X"1A",X"00",X"F7",X"57",X"01",X"00",
		X"21",X"03",X"4E",X"34",X"C9",X"21",X"15",X"4E",X"35",X"CD",X"E4",X"29",X"AF",X"32",X"79",X"4C",
		X"AF",X"32",X"03",X"4E",X"32",X"02",X"4E",X"32",X"04",X"4E",X"21",X"00",X"4E",X"34",X"C9",X"3A",
		X"04",X"4E",X"E7",X"D6",X"0A",X"F6",X"0A",X"0C",X"00",X"2A",X"0B",X"6D",X"0B",X"0C",X"00",X"BA",
		X"0B",X"0C",X"00",X"05",X"0C",X"22",X"0C",X"0C",X"00",X"75",X"0C",X"7B",X"0C",X"0C",X"00",X"8B",
		X"0C",X"0C",X"00",X"A1",X"0C",X"0C",X"00",X"A5",X"0C",X"0C",X"00",X"A7",X"0C",X"0C",X"00",X"A9",
		X"0C",X"0C",X"00",X"AB",X"0C",X"0C",X"00",X"AD",X"0C",X"0C",X"00",X"AF",X"0C",X"0C",X"00",X"B1",
		X"0C",X"0C",X"00",X"CF",X"0C",X"0C",X"00",X"17",X"0D",X"3B",X"0D",X"0C",X"00",X"3E",X"0D",X"0C",
		X"00",X"84",X"B1",X"5F",X"09",X"5F",X"09",X"5F",X"09",X"A6",X"3F",X"0C",X"00",X"A9",X"68",X"0C",
		X"00",X"54",X"76",X"0C",X"00",X"E0",X"7F",X"0C",X"00",X"E0",X"7F",X"0C",X"00",X"E0",X"7F",X"3E",
		X"27",X"32",X"04",X"4E",X"C9",X"78",X"A7",X"20",X"04",X"2A",X"0A",X"4E",X"7E",X"DD",X"21",X"ED",
		X"09",X"47",X"87",X"87",X"80",X"80",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"7E",X"00",X"87",X"47",
		X"87",X"87",X"4F",X"87",X"87",X"81",X"80",X"5F",X"16",X"00",X"21",X"A5",X"32",X"19",X"CD",X"6B",
		X"0A",X"DD",X"7E",X"01",X"32",X"B0",X"4D",X"DD",X"7E",X"02",X"47",X"87",X"80",X"5F",X"16",X"00",
		X"21",X"9A",X"0A",X"19",X"CD",X"91",X"0A",X"DD",X"7E",X"03",X"87",X"5F",X"16",X"00",X"FD",X"21",
		X"A6",X"0A",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"22",X"BB",X"4D",X"DD",X"7E",X"04",
		X"87",X"5F",X"16",X"00",X"FD",X"21",X"B8",X"0A",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",
		X"22",X"BD",X"4D",X"DD",X"7E",X"05",X"87",X"5F",X"16",X"00",X"FD",X"21",X"D0",X"0A",X"FD",X"19",
		X"FD",X"6E",X"00",X"FD",X"66",X"01",X"22",X"95",X"4D",X"CD",X"64",X"2A",X"C9",X"03",X"01",X"01",
		X"00",X"02",X"00",X"04",X"01",X"02",X"01",X"03",X"00",X"04",X"01",X"03",X"02",X"04",X"01",X"04",
		X"02",X"03",X"02",X"05",X"01",X"05",X"00",X"03",X"02",X"06",X"02",X"05",X"01",X"03",X"03",X"03",
		X"02",X"05",X"02",X"03",X"03",X"06",X"02",X"05",X"02",X"03",X"03",X"06",X"02",X"05",X"00",X"03",
		X"04",X"07",X"02",X"05",X"01",X"03",X"04",X"03",X"02",X"05",X"02",X"03",X"04",X"06",X"02",X"05",
		X"02",X"03",X"05",X"07",X"02",X"05",X"00",X"03",X"05",X"07",X"02",X"05",X"02",X"03",X"05",X"05",
		X"02",X"05",X"01",X"03",X"06",X"07",X"02",X"05",X"02",X"03",X"06",X"07",X"02",X"05",X"02",X"03",
		X"06",X"08",X"02",X"05",X"02",X"03",X"06",X"07",X"02",X"05",X"02",X"03",X"07",X"08",X"02",X"05",
		X"02",X"03",X"07",X"08",X"02",X"06",X"02",X"03",X"07",X"08",X"02",X"11",X"46",X"4D",X"01",X"1C",
		X"00",X"ED",X"B0",X"01",X"0C",X"00",X"A7",X"ED",X"42",X"ED",X"B0",X"01",X"0C",X"00",X"A7",X"ED",
		X"42",X"ED",X"B0",X"01",X"0C",X"00",X"A7",X"ED",X"42",X"ED",X"B0",X"01",X"0E",X"00",X"ED",X"B0",
		X"C9",X"11",X"B8",X"4D",X"01",X"03",X"00",X"ED",X"B0",X"C9",X"14",X"1E",X"46",X"00",X"1E",X"3C",
		X"00",X"00",X"32",X"00",X"00",X"00",X"14",X"0A",X"1E",X"0F",X"28",X"14",X"32",X"19",X"3C",X"1E",
		X"50",X"28",X"64",X"32",X"78",X"3C",X"8C",X"46",X"C0",X"03",X"48",X"03",X"D0",X"02",X"58",X"02",
		X"E0",X"01",X"E0",X"01",X"68",X"01",X"68",X"01",X"F0",X"00",X"F0",X"00",X"78",X"00",X"01",X"00",
		X"F0",X"00",X"F0",X"00",X"B4",X"00",X"21",X"09",X"4E",X"AF",X"06",X"0B",X"CF",X"CD",X"B5",X"22",
		X"2A",X"73",X"4E",X"22",X"0A",X"4E",X"21",X"0A",X"4E",X"11",X"38",X"4E",X"01",X"2E",X"00",X"ED",
		X"B0",X"21",X"04",X"4E",X"34",X"C9",X"3A",X"00",X"4E",X"3D",X"20",X"06",X"3E",X"09",X"32",X"04",
		X"4E",X"C9",X"EF",X"11",X"00",X"EF",X"1C",X"83",X"EF",X"04",X"00",X"EF",X"05",X"00",X"EF",X"10",
		X"00",X"EF",X"1A",X"00",X"F7",X"54",X"00",X"00",X"F7",X"54",X"06",X"00",X"3A",X"72",X"4E",X"47",
		X"3A",X"09",X"4E",X"A0",X"32",X"03",X"50",X"C3",X"F1",X"0A",X"3A",X"00",X"50",X"CB",X"67",X"C3",
		X"3B",X"0B",X"21",X"04",X"4E",X"36",X"0E",X"EF",X"13",X"00",X"C9",X"3A",X"0E",X"4E",X"C3",X"7A",
		X"94",X"00",X"21",X"04",X"4E",X"36",X"0C",X"C9",X"CD",X"B7",X"11",X"CD",X"B7",X"11",X"CD",X"14",
		X"16",X"CD",X"1F",X"0F",X"CD",X"00",X"11",X"CD",X"19",X"11",X"CD",X"5E",X"0D",X"CD",X"BC",X"0E",
		X"CD",X"F3",X"0E",X"CD",X"FA",X"B2",X"CD",X"4E",X"11",X"CD",X"8F",X"11",X"C9",X"3E",X"01",X"32",
		X"12",X"4E",X"CD",X"8A",X"22",X"21",X"04",X"4E",X"34",X"3A",X"14",X"4E",X"A7",X"20",X"39",X"3A",
		X"70",X"4E",X"A7",X"28",X"33",X"3A",X"42",X"4E",X"A7",X"28",X"2D",X"3A",X"09",X"4E",X"C6",X"03",
		X"4F",X"06",X"1C",X"CD",X"42",X"00",X"EF",X"1C",X"05",X"3A",X"FE",X"4D",X"A7",X"20",X"05",X"F7",
		X"54",X"00",X"00",X"C9",X"3D",X"47",X"3A",X"09",X"4E",X"B8",X"C0",X"3A",X"04",X"4E",X"3C",X"32",
		X"FF",X"4D",X"3E",X"27",X"32",X"04",X"4E",X"C9",X"34",X"C9",X"3A",X"70",X"4E",X"A7",X"28",X"06",
		X"3A",X"42",X"4E",X"A7",X"20",X"2E",X"3A",X"14",X"4E",X"A7",X"20",X"33",X"CD",X"1B",X"2A",X"EF",
		X"1C",X"05",X"3A",X"FE",X"4D",X"A7",X"20",X"06",X"F7",X"54",X"00",X"00",X"18",X"11",X"21",X"04",
		X"4E",X"34",X"34",X"3A",X"04",X"4E",X"32",X"FF",X"4D",X"3E",X"27",X"32",X"04",X"4E",X"C9",X"21",
		X"04",X"4E",X"34",X"C9",X"CD",X"41",X"0D",X"3A",X"09",X"4E",X"EE",X"01",X"32",X"09",X"4E",X"3E",
		X"09",X"32",X"04",X"4E",X"C9",X"3A",X"78",X"4C",X"3C",X"32",X"78",X"4C",X"AF",X"32",X"02",X"4E",
		X"32",X"04",X"4E",X"32",X"70",X"4E",X"32",X"09",X"4E",X"32",X"03",X"50",X"3E",X"01",X"32",X"00",
		X"4E",X"C9",X"EF",X"00",X"01",X"EF",X"01",X"01",X"EF",X"02",X"00",X"EF",X"11",X"00",X"EF",X"13",
		X"00",X"EF",X"03",X"00",X"EF",X"04",X"00",X"EF",X"05",X"00",X"EF",X"1C",X"0E",X"EF",X"10",X"00",
		X"EF",X"1A",X"00",X"EF",X"1C",X"06",X"EF",X"29",X"0F",X"EF",X"37",X"0F",X"3A",X"00",X"4E",X"FE",
		X"03",X"28",X"06",X"EF",X"1C",X"05",X"EF",X"1D",X"00",X"F7",X"54",X"00",X"00",X"3A",X"00",X"4E",
		X"3D",X"28",X"04",X"F7",X"54",X"06",X"00",X"3A",X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"32",
		X"03",X"50",X"C3",X"F1",X"0A",X"3E",X"03",X"32",X"04",X"4E",X"C9",X"F7",X"54",X"00",X"00",X"21",
		X"04",X"4E",X"34",X"AF",X"32",X"AC",X"4E",X"32",X"BC",X"4E",X"C9",X"0E",X"02",X"06",X"01",X"CD",
		X"42",X"00",X"F7",X"42",X"00",X"00",X"21",X"00",X"00",X"CD",X"68",X"24",X"21",X"04",X"4E",X"34",
		X"C9",X"0E",X"00",X"18",X"E8",X"18",X"E4",X"18",X"F8",X"18",X"E0",X"18",X"F4",X"18",X"DC",X"18",
		X"F0",X"EF",X"00",X"01",X"EF",X"06",X"00",X"EF",X"11",X"00",X"EF",X"13",X"00",X"EF",X"04",X"01",
		X"EF",X"05",X"01",X"EF",X"10",X"13",X"F7",X"43",X"00",X"00",X"21",X"04",X"4E",X"34",X"C9",X"AF",
		X"32",X"AC",X"4E",X"32",X"BC",X"4E",X"3A",X"13",X"4E",X"FE",X"14",X"38",X"02",X"3E",X"14",X"E7",
		X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",
		X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",
		X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"0A",X"0D",X"21",X"04",X"4E",X"34",X"34",X"AF",
		X"32",X"CC",X"4E",X"32",X"DC",X"4E",X"C9",X"AF",X"32",X"CC",X"4E",X"32",X"DC",X"4E",X"06",X"07",
		X"21",X"0C",X"4E",X"CF",X"CD",X"B5",X"22",X"21",X"04",X"4E",X"34",X"21",X"13",X"4E",X"34",X"2A",
		X"0A",X"4E",X"7E",X"FE",X"14",X"C8",X"23",X"22",X"0A",X"4E",X"C9",X"C3",X"22",X"0C",X"C3",X"75",
		X"0C",X"06",X"2E",X"DD",X"21",X"0A",X"4E",X"FD",X"21",X"38",X"4E",X"DD",X"56",X"00",X"FD",X"5E",
		X"00",X"FD",X"72",X"00",X"DD",X"73",X"00",X"DD",X"23",X"FD",X"23",X"10",X"EE",X"C9",X"3A",X"A4",
		X"4D",X"A7",X"C0",X"DD",X"21",X"00",X"4C",X"FD",X"21",X"C8",X"4D",X"11",X"00",X"01",X"FD",X"BE",
		X"00",X"C2",X"B8",X"0E",X"FD",X"36",X"00",X"0E",X"3A",X"A6",X"4D",X"A7",X"28",X"26",X"2A",X"CB",
		X"4D",X"A7",X"ED",X"52",X"30",X"1E",X"21",X"AC",X"4E",X"CB",X"FE",X"3E",X"09",X"DD",X"BE",X"0B",
		X"20",X"02",X"CB",X"BE",X"3A",X"D2",X"4F",X"CB",X"47",X"28",X"04",X"3E",X"05",X"18",X"02",X"3E",
		X"09",X"32",X"0B",X"4C",X"3A",X"A7",X"4D",X"A7",X"28",X"2D",X"2A",X"CB",X"4D",X"A7",X"ED",X"52",
		X"30",X"37",X"3E",X"11",X"DD",X"BE",X"03",X"28",X"0F",X"3A",X"70",X"4C",X"FE",X"03",X"CA",X"E9",
		X"0D",X"DD",X"36",X"03",X"11",X"C3",X"E9",X"0D",X"3A",X"70",X"4C",X"FE",X"03",X"CA",X"E9",X"0D",
		X"DD",X"36",X"03",X"12",X"C3",X"E9",X"0D",X"3E",X"01",X"DD",X"BE",X"03",X"28",X"07",X"DD",X"36",
		X"03",X"01",X"C3",X"E9",X"0D",X"DD",X"36",X"03",X"01",X"3A",X"A8",X"4D",X"A7",X"28",X"2D",X"2A",
		X"CB",X"4D",X"A7",X"ED",X"52",X"30",X"37",X"3E",X"11",X"DD",X"BE",X"05",X"28",X"0F",X"3A",X"70",
		X"4C",X"FE",X"03",X"CA",X"2E",X"0E",X"DD",X"36",X"05",X"11",X"C3",X"2E",X"0E",X"3A",X"70",X"4C",
		X"FE",X"03",X"CA",X"2E",X"0E",X"DD",X"36",X"05",X"12",X"C3",X"2E",X"0E",X"3E",X"03",X"DD",X"BE",
		X"05",X"28",X"07",X"DD",X"36",X"05",X"03",X"C3",X"2E",X"0E",X"DD",X"36",X"05",X"03",X"3A",X"A9",
		X"4D",X"A7",X"28",X"2D",X"2A",X"CB",X"4D",X"A7",X"ED",X"52",X"30",X"37",X"3E",X"11",X"DD",X"BE",
		X"07",X"28",X"0F",X"3A",X"70",X"4C",X"FE",X"03",X"CA",X"73",X"0E",X"DD",X"36",X"07",X"11",X"C3",
		X"73",X"0E",X"3A",X"70",X"4C",X"FE",X"03",X"CA",X"73",X"0E",X"DD",X"36",X"07",X"12",X"C3",X"73",
		X"0E",X"3E",X"05",X"DD",X"BE",X"07",X"28",X"07",X"DD",X"36",X"07",X"05",X"C3",X"73",X"0E",X"DD",
		X"36",X"07",X"05",X"3A",X"AA",X"4D",X"A7",X"28",X"2D",X"2A",X"CB",X"4D",X"A7",X"ED",X"52",X"30",
		X"37",X"3E",X"11",X"DD",X"BE",X"09",X"28",X"0F",X"3A",X"70",X"4C",X"FE",X"03",X"CA",X"B8",X"0E",
		X"DD",X"36",X"09",X"11",X"C3",X"B8",X"0E",X"3A",X"70",X"4C",X"FE",X"03",X"CA",X"B8",X"0E",X"DD",
		X"36",X"09",X"12",X"C3",X"B8",X"0E",X"3E",X"07",X"DD",X"BE",X"09",X"28",X"07",X"DD",X"36",X"09",
		X"07",X"C3",X"B8",X"0E",X"DD",X"36",X"09",X"07",X"FD",X"35",X"00",X"C9",X"06",X"19",X"3A",X"02",
		X"4E",X"FE",X"27",X"C2",X"C8",X"0E",X"06",X"00",X"DD",X"21",X"00",X"4C",X"3A",X"AC",X"4D",X"A7",
		X"CA",X"D6",X"0E",X"DD",X"70",X"03",X"3A",X"AD",X"4D",X"A7",X"CA",X"E0",X"0E",X"DD",X"70",X"05",
		X"3A",X"AE",X"4D",X"A7",X"CA",X"EA",X"0E",X"DD",X"70",X"07",X"3A",X"AF",X"4D",X"A7",X"C8",X"DD",
		X"70",X"09",X"C9",X"3A",X"70",X"4C",X"FE",X"03",X"C8",X"21",X"CF",X"4D",X"34",X"3E",X"0A",X"BE",
		X"C0",X"36",X"00",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"06",X"21",X"64",X"44",X"C3",X"3D",X"95",
		X"21",X"32",X"47",X"3E",X"10",X"BE",X"20",X"02",X"3E",X"00",X"77",X"32",X"78",X"46",X"C9",X"3A",
		X"A4",X"4D",X"A7",X"C0",X"3A",X"94",X"4D",X"07",X"32",X"94",X"4D",X"D0",X"3A",X"A0",X"4D",X"A7",
		X"C2",X"6D",X"0F",X"DD",X"21",X"8B",X"32",X"FD",X"21",X"00",X"4D",X"CD",X"CD",X"1E",X"22",X"00",
		X"4D",X"3E",X"03",X"32",X"28",X"4D",X"32",X"2C",X"4D",X"3A",X"00",X"4D",X"FE",X"64",X"C2",X"6D",
		X"0F",X"21",X"2C",X"2E",X"22",X"0A",X"4D",X"21",X"00",X"01",X"22",X"14",X"4D",X"22",X"1E",X"4D",
		X"3E",X"02",X"32",X"28",X"4D",X"32",X"2C",X"4D",X"3E",X"01",X"32",X"A0",X"4D",X"3A",X"A1",X"4D",
		X"FE",X"01",X"CA",X"D8",X"0F",X"FE",X"00",X"C2",X"9E",X"0F",X"3A",X"02",X"4D",X"FE",X"78",X"CC",
		X"AD",X"2E",X"FE",X"80",X"CC",X"AD",X"2E",X"3A",X"2D",X"4D",X"32",X"29",X"4D",X"DD",X"21",X"20",
		X"4D",X"FD",X"21",X"02",X"4D",X"CD",X"CD",X"1E",X"22",X"02",X"4D",X"C3",X"D8",X"0F",X"DD",X"21",
		X"8B",X"32",X"FD",X"21",X"02",X"4D",X"CD",X"CD",X"1E",X"22",X"02",X"4D",X"3E",X"03",X"32",X"2D",
		X"4D",X"32",X"29",X"4D",X"3A",X"02",X"4D",X"FE",X"64",X"C2",X"D8",X"0F",X"21",X"2C",X"2E",X"22",
		X"0C",X"4D",X"21",X"00",X"01",X"22",X"16",X"4D",X"22",X"20",X"4D",X"3E",X"02",X"32",X"29",X"4D",
		X"32",X"2D",X"4D",X"3E",X"01",X"32",X"A1",X"4D",X"3A",X"A2",X"4D",X"FE",X"01",X"CA",X"70",X"10",
		X"FE",X"00",X"C2",X"09",X"10",X"3A",X"04",X"4D",X"FE",X"78",X"CC",X"D4",X"2E",X"FE",X"80",X"CC",
		X"D4",X"2E",X"3A",X"2E",X"4D",X"32",X"2A",X"4D",X"DD",X"21",X"22",X"4D",X"FD",X"21",X"04",X"4D",
		X"CD",X"CD",X"1E",X"22",X"04",X"4D",X"C3",X"70",X"10",X"3A",X"A2",X"4D",X"FE",X"03",X"C2",X"36",
		X"10",X"DD",X"21",X"85",X"32",X"FD",X"21",X"04",X"4D",X"CD",X"CD",X"1E",X"22",X"04",X"4D",X"AF",
		X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"3A",X"05",X"4D",X"FE",X"80",X"C2",X"70",X"10",X"3E",X"02",
		X"32",X"A2",X"4D",X"C3",X"70",X"10",X"DD",X"21",X"8B",X"32",X"FD",X"21",X"04",X"4D",X"CD",X"CD",
		X"1E",X"22",X"04",X"4D",X"3E",X"03",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"3A",X"04",X"4D",X"FE",
		X"64",X"C2",X"70",X"10",X"21",X"2C",X"2E",X"22",X"0E",X"4D",X"21",X"00",X"01",X"22",X"18",X"4D",
		X"22",X"22",X"4D",X"3E",X"02",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"3E",X"01",X"32",X"A2",X"4D",
		X"3A",X"A3",X"4D",X"FE",X"01",X"C8",X"FE",X"00",X"C2",X"9D",X"10",X"3A",X"06",X"4D",X"FE",X"78",
		X"CC",X"FB",X"2E",X"FE",X"80",X"CC",X"FB",X"2E",X"3A",X"2F",X"4D",X"32",X"2B",X"4D",X"DD",X"21",
		X"24",X"4D",X"FD",X"21",X"06",X"4D",X"CD",X"CD",X"1E",X"22",X"06",X"4D",X"C9",X"3A",X"A3",X"4D",
		X"FE",X"03",X"C2",X"C7",X"10",X"DD",X"21",X"89",X"32",X"FD",X"21",X"06",X"4D",X"CD",X"CD",X"1E",
		X"22",X"06",X"4D",X"3E",X"02",X"32",X"2B",X"4D",X"32",X"2F",X"4D",X"3A",X"07",X"4D",X"FE",X"80",
		X"C0",X"3E",X"02",X"32",X"A3",X"4D",X"C9",X"DD",X"21",X"8B",X"32",X"FD",X"21",X"06",X"4D",X"CD",
		X"CD",X"1E",X"22",X"06",X"4D",X"3E",X"03",X"32",X"2B",X"4D",X"32",X"2F",X"4D",X"3A",X"06",X"4D",
		X"FE",X"64",X"C0",X"21",X"2C",X"2E",X"22",X"10",X"4D",X"21",X"00",X"01",X"22",X"1A",X"4D",X"22",
		X"24",X"4D",X"3E",X"02",X"32",X"2B",X"4D",X"32",X"2F",X"4D",X"3E",X"01",X"32",X"A3",X"4D",X"C9",
		X"21",X"C4",X"4D",X"34",X"3E",X"08",X"BE",X"C0",X"36",X"00",X"3A",X"70",X"4C",X"FE",X"03",X"C8",
		X"3A",X"C0",X"4D",X"EE",X"01",X"32",X"C0",X"4D",X"C9",X"3A",X"A6",X"4D",X"A7",X"C0",X"3A",X"C1",
		X"4D",X"FE",X"07",X"C8",X"87",X"2A",X"C2",X"4D",X"23",X"22",X"C2",X"4D",X"5F",X"16",X"00",X"DD",
		X"21",X"86",X"4D",X"DD",X"19",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"A7",X"ED",X"52",X"C0",X"AF",
		X"3C",X"32",X"C1",X"4D",X"21",X"01",X"01",X"22",X"B1",X"4D",X"22",X"B3",X"4D",X"C9",X"3A",X"A5",
		X"4D",X"A7",X"28",X"05",X"AF",X"32",X"AC",X"4E",X"C9",X"21",X"AC",X"4E",X"06",X"E0",X"3A",X"0E",
		X"4E",X"FE",X"E4",X"38",X"06",X"78",X"A6",X"CB",X"E7",X"77",X"C9",X"FE",X"D4",X"38",X"06",X"78",
		X"A6",X"CB",X"DF",X"77",X"C9",X"FE",X"B4",X"38",X"06",X"78",X"A6",X"CB",X"D7",X"77",X"C9",X"FE",
		X"74",X"38",X"06",X"78",X"A6",X"CB",X"CF",X"77",X"C9",X"78",X"A6",X"CB",X"C7",X"77",X"C9",X"3A",
		X"70",X"4C",X"FE",X"03",X"C8",X"FE",X"02",X"CC",X"79",X"85",X"CD",X"A0",X"11",X"C3",X"79",X"85",
		X"3A",X"0E",X"4E",X"FE",X"A0",X"D8",X"3A",X"70",X"4C",X"FE",X"02",X"CC",X"79",X"85",X"C9",X"AF",
		X"32",X"D4",X"4D",X"C9",X"C3",X"D7",X"35",X"CD",X"B1",X"14",X"3A",X"A5",X"4D",X"A7",X"C0",X"CD",
		X"58",X"12",X"CD",X"86",X"12",X"CD",X"96",X"12",X"CD",X"A6",X"12",X"CD",X"B8",X"12",X"3A",X"A4",
		X"4D",X"A7",X"CA",X"D9",X"11",X"CD",X"3F",X"14",X"C9",X"CD",X"96",X"19",X"CD",X"02",X"1A",X"3A",
		X"A4",X"4D",X"A7",X"C0",X"CD",X"7F",X"1A",X"3A",X"70",X"4C",X"A7",X"28",X"27",X"3A",X"70",X"4C",
		X"FE",X"01",X"28",X"20",X"3A",X"72",X"4C",X"A7",X"28",X"1A",X"CD",X"7F",X"1A",X"CD",X"2E",X"A3",
		X"3A",X"13",X"4E",X"FE",X"05",X"38",X"0D",X"CD",X"F1",X"A5",X"3A",X"13",X"4E",X"FE",X"10",X"38",
		X"03",X"CD",X"1A",X"A5",X"CD",X"2E",X"A3",X"CD",X"43",X"A4",X"CD",X"1A",X"A5",X"CD",X"F1",X"A5",
		X"3A",X"13",X"4E",X"FE",X"08",X"38",X"1E",X"CD",X"F1",X"A5",X"3A",X"70",X"4C",X"FE",X"03",X"20",
		X"14",X"3A",X"13",X"4E",X"FE",X"0B",X"38",X"0D",X"CD",X"1A",X"A5",X"3A",X"0E",X"4E",X"FE",X"A0",
		X"38",X"03",X"CD",X"2E",X"A3",X"3A",X"04",X"4E",X"FE",X"03",X"C0",X"CD",X"A2",X"15",X"CD",X"33",
		X"1F",X"CD",X"56",X"1F",X"CD",X"79",X"1F",X"C9",X"3A",X"AB",X"4D",X"A7",X"C8",X"3D",X"20",X"08",
		X"32",X"AB",X"4D",X"3C",X"32",X"AC",X"4D",X"C9",X"3D",X"20",X"08",X"32",X"AB",X"4D",X"3C",X"32",
		X"AD",X"4D",X"C9",X"3D",X"20",X"08",X"32",X"AB",X"4D",X"3C",X"32",X"AE",X"4D",X"C9",X"32",X"AF",
		X"4D",X"3D",X"32",X"AB",X"4D",X"C9",X"3A",X"AC",X"4D",X"E6",X"03",X"E7",X"0C",X"00",X"CA",X"12",
		X"DC",X"12",X"80",X"67",X"90",X"68",X"3A",X"AD",X"4D",X"E6",X"03",X"E7",X"0C",X"00",X"22",X"13",
		X"34",X"13",X"80",X"67",X"90",X"68",X"3A",X"AE",X"4D",X"E6",X"03",X"E7",X"0C",X"00",X"66",X"13",
		X"78",X"13",X"99",X"13",X"00",X"60",X"00",X"67",X"3A",X"AF",X"4D",X"E6",X"03",X"E7",X"0C",X"00",
		X"D3",X"13",X"E5",X"13",X"06",X"14",X"A0",X"67",X"A0",X"67",X"CD",X"D0",X"A3",X"2A",X"00",X"4D",
		X"11",X"64",X"80",X"A7",X"ED",X"52",X"C0",X"21",X"AC",X"4D",X"34",X"C9",X"DD",X"21",X"87",X"32",
		X"FD",X"21",X"00",X"4D",X"CD",X"CD",X"1E",X"22",X"00",X"4D",X"3E",X"01",X"32",X"28",X"4D",X"32",
		X"2C",X"4D",X"3A",X"00",X"4D",X"FE",X"80",X"C0",X"21",X"2F",X"2E",X"22",X"0A",X"4D",X"22",X"31",
		X"4D",X"AF",X"32",X"A0",X"4D",X"32",X"AC",X"4D",X"32",X"A7",X"4D",X"DD",X"21",X"AC",X"4D",X"DD",
		X"B6",X"00",X"DD",X"B6",X"01",X"DD",X"B6",X"02",X"DD",X"B6",X"03",X"C0",X"21",X"AC",X"4E",X"CB",
		X"B6",X"C9",X"CD",X"A7",X"A4",X"2A",X"02",X"4D",X"11",X"64",X"80",X"A7",X"ED",X"52",X"C0",X"21",
		X"AD",X"4D",X"34",X"C9",X"DD",X"21",X"87",X"32",X"FD",X"21",X"02",X"4D",X"CD",X"CD",X"1E",X"22",
		X"02",X"4D",X"3E",X"01",X"32",X"29",X"4D",X"32",X"2D",X"4D",X"3A",X"02",X"4D",X"FE",X"80",X"C0",
		X"21",X"2F",X"2E",X"22",X"0C",X"4D",X"22",X"33",X"4D",X"AF",X"32",X"A1",X"4D",X"32",X"AD",X"4D",
		X"32",X"A8",X"4D",X"C3",X"0B",X"13",X"CD",X"7E",X"A5",X"2A",X"04",X"4D",X"11",X"64",X"80",X"A7",
		X"ED",X"52",X"C0",X"21",X"AE",X"4D",X"34",X"C9",X"DD",X"21",X"87",X"32",X"FD",X"21",X"04",X"4D",
		X"CD",X"CD",X"1E",X"22",X"04",X"4D",X"3E",X"01",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"3A",X"04",
		X"4D",X"FE",X"80",X"C0",X"21",X"AE",X"4D",X"34",X"C9",X"DD",X"21",X"89",X"32",X"FD",X"21",X"04",
		X"4D",X"CD",X"CD",X"1E",X"22",X"04",X"4D",X"3E",X"02",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"3A",
		X"05",X"4D",X"FE",X"90",X"C0",X"21",X"2F",X"30",X"22",X"0E",X"4D",X"22",X"35",X"4D",X"3E",X"01",
		X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"AF",X"32",X"A2",X"4D",X"32",X"AE",X"4D",X"32",X"A9",X"4D",
		X"C3",X"0B",X"13",X"CD",X"55",X"A6",X"2A",X"06",X"4D",X"11",X"64",X"80",X"A7",X"ED",X"52",X"C0",
		X"21",X"AF",X"4D",X"34",X"C9",X"DD",X"21",X"87",X"32",X"FD",X"21",X"06",X"4D",X"CD",X"CD",X"1E",
		X"22",X"06",X"4D",X"3E",X"01",X"32",X"2B",X"4D",X"32",X"2F",X"4D",X"3A",X"06",X"4D",X"FE",X"80",
		X"C0",X"21",X"AF",X"4D",X"34",X"C9",X"DD",X"21",X"85",X"32",X"FD",X"21",X"06",X"4D",X"CD",X"CD",
		X"1E",X"22",X"06",X"4D",X"AF",X"32",X"2B",X"4D",X"32",X"2F",X"4D",X"3A",X"07",X"4D",X"FE",X"70",
		X"C0",X"21",X"2F",X"2C",X"22",X"10",X"4D",X"22",X"37",X"4D",X"3E",X"01",X"32",X"2B",X"4D",X"32",
		X"2F",X"4D",X"AF",X"32",X"A3",X"4D",X"32",X"AF",X"4D",X"32",X"AA",X"4D",X"C3",X"0B",X"13",X"3A",
		X"D1",X"4D",X"E6",X"03",X"E7",X"4D",X"14",X"0C",X"00",X"4D",X"14",X"0C",X"00",X"21",X"00",X"4C",
		X"3A",X"A4",X"4D",X"87",X"5F",X"16",X"00",X"19",X"3A",X"D1",X"4D",X"A7",X"20",X"2E",X"3A",X"D0",
		X"4D",X"06",X"27",X"80",X"47",X"3A",X"72",X"4E",X"4F",X"3A",X"09",X"4E",X"A1",X"28",X"04",X"CB",
		X"F0",X"CB",X"F8",X"70",X"23",X"36",X"18",X"3A",X"70",X"4C",X"FE",X"03",X"28",X"02",X"3E",X"00",
		X"32",X"0B",X"4C",X"F7",X"4A",X"03",X"00",X"21",X"D1",X"4D",X"34",X"C9",X"36",X"20",X"3A",X"D2",
		X"4F",X"CB",X"47",X"20",X"04",X"3E",X"09",X"18",X"02",X"3E",X"05",X"32",X"0B",X"4C",X"3A",X"A4",
		X"4D",X"32",X"AB",X"4D",X"AF",X"32",X"A4",X"4D",X"32",X"D1",X"4D",X"21",X"AC",X"4E",X"CB",X"F6",
		X"C9",X"3A",X"A5",X"4D",X"E7",X"0C",X"00",X"E3",X"14",X"E3",X"14",X"E3",X"14",X"E3",X"14",X"F7",
		X"14",X"25",X"15",X"32",X"15",X"3A",X"15",X"42",X"15",X"4A",X"15",X"52",X"15",X"5A",X"15",X"62",
		X"15",X"6A",X"15",X"72",X"15",X"7F",X"15",X"50",X"65",X"50",X"65",X"80",X"67",X"80",X"67",X"50",
		X"65",X"80",X"67",X"2A",X"C5",X"4D",X"23",X"22",X"C5",X"4D",X"11",X"78",X"00",X"A7",X"ED",X"52",
		X"C0",X"3E",X"05",X"32",X"A5",X"4D",X"C9",X"21",X"00",X"00",X"CD",X"68",X"24",X"3E",X"34",X"11",
		X"B4",X"00",X"4F",X"3A",X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"28",X"04",X"3E",X"C0",X"B1",
		X"4F",X"79",X"32",X"0A",X"4C",X"2A",X"C5",X"4D",X"23",X"22",X"C5",X"4D",X"A7",X"ED",X"52",X"C0",
		X"21",X"A5",X"4D",X"34",X"C9",X"21",X"BC",X"4E",X"CB",X"E6",X"3E",X"35",X"11",X"C3",X"00",X"C3",
		X"02",X"15",X"3E",X"36",X"11",X"D2",X"00",X"C3",X"02",X"15",X"3E",X"37",X"11",X"E1",X"00",X"C3",
		X"02",X"15",X"3E",X"38",X"11",X"F0",X"00",X"C3",X"02",X"15",X"3E",X"39",X"11",X"FF",X"00",X"C3",
		X"02",X"15",X"3E",X"3A",X"11",X"0E",X"01",X"C3",X"02",X"15",X"3E",X"3B",X"11",X"1D",X"01",X"C3",
		X"02",X"15",X"3E",X"3C",X"11",X"2C",X"01",X"C3",X"02",X"15",X"3E",X"3D",X"11",X"3B",X"01",X"C3",
		X"02",X"15",X"21",X"BC",X"4E",X"36",X"00",X"3E",X"3E",X"11",X"59",X"01",X"C3",X"02",X"15",X"3E",
		X"3F",X"32",X"0A",X"4C",X"2A",X"C5",X"4D",X"23",X"22",X"C5",X"4D",X"11",X"B8",X"01",X"A7",X"ED",
		X"52",X"C0",X"21",X"14",X"4E",X"35",X"21",X"15",X"4E",X"35",X"CD",X"5F",X"24",X"21",X"04",X"4E",
		X"34",X"C9",X"3A",X"A6",X"4D",X"A7",X"C8",X"DD",X"21",X"A7",X"4D",X"DD",X"7E",X"00",X"DD",X"B6",
		X"01",X"DD",X"B6",X"02",X"DD",X"B6",X"03",X"CA",X"C4",X"15",X"2A",X"CB",X"4D",X"2B",X"22",X"CB",
		X"4D",X"7C",X"B5",X"C0",X"21",X"0B",X"4C",X"3A",X"D2",X"4F",X"CB",X"47",X"20",X"04",X"36",X"09",
		X"18",X"02",X"36",X"05",X"3A",X"AC",X"4D",X"A7",X"C2",X"DE",X"15",X"32",X"A7",X"4D",X"3A",X"AD",
		X"4D",X"A7",X"C2",X"E8",X"15",X"32",X"A8",X"4D",X"3A",X"AE",X"4D",X"A7",X"C2",X"F2",X"15",X"32",
		X"A9",X"4D",X"3A",X"AF",X"4D",X"A7",X"C2",X"FC",X"15",X"32",X"AA",X"4D",X"AF",X"32",X"CB",X"4D",
		X"32",X"CC",X"4D",X"32",X"A6",X"4D",X"32",X"C8",X"4D",X"32",X"D0",X"4D",X"21",X"AC",X"4E",X"CB",
		X"AE",X"CB",X"BE",X"C9",X"21",X"9E",X"4D",X"3A",X"0E",X"4E",X"BE",X"CA",X"25",X"16",X"21",X"00",
		X"00",X"22",X"97",X"4D",X"C9",X"2A",X"97",X"4D",X"23",X"22",X"97",X"4D",X"ED",X"5B",X"95",X"4D",
		X"A7",X"ED",X"52",X"C0",X"21",X"00",X"00",X"22",X"97",X"4D",X"3A",X"A1",X"4D",X"A7",X"F5",X"CC",
		X"50",X"1F",X"F1",X"C8",X"3A",X"A2",X"4D",X"A7",X"F5",X"CC",X"73",X"1F",X"F1",X"C8",X"3A",X"A3",
		X"4D",X"A7",X"CC",X"9B",X"1F",X"C9",X"3A",X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"C8",X"47",
		X"DD",X"21",X"00",X"4C",X"1E",X"08",X"0E",X"08",X"16",X"07",X"3A",X"00",X"4D",X"83",X"DD",X"77",
		X"13",X"3A",X"01",X"4D",X"2F",X"82",X"DD",X"77",X"12",X"3A",X"02",X"4D",X"83",X"DD",X"77",X"15",
		X"3A",X"03",X"4D",X"2F",X"82",X"DD",X"77",X"14",X"3A",X"04",X"4D",X"83",X"DD",X"77",X"17",X"3A",
		X"05",X"4D",X"2F",X"81",X"DD",X"77",X"16",X"3A",X"06",X"4D",X"83",X"DD",X"77",X"19",X"3A",X"07",
		X"4D",X"2F",X"81",X"DD",X"77",X"18",X"3A",X"08",X"4D",X"83",X"DD",X"77",X"1B",X"3A",X"09",X"4D",
		X"2F",X"81",X"DD",X"77",X"1A",X"3A",X"D2",X"4D",X"83",X"DD",X"77",X"1D",X"3A",X"D3",X"4D",X"2F",
		X"81",X"DD",X"77",X"1C",X"C3",X"35",X"17",X"3A",X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"C0",
		X"47",X"1E",X"09",X"0E",X"07",X"16",X"06",X"DD",X"21",X"00",X"4C",X"3A",X"00",X"4D",X"2F",X"83",
		X"DD",X"77",X"13",X"3A",X"01",X"4D",X"82",X"DD",X"77",X"12",X"3A",X"02",X"4D",X"2F",X"83",X"DD",
		X"77",X"15",X"3A",X"03",X"4D",X"82",X"DD",X"77",X"14",X"3A",X"04",X"4D",X"2F",X"83",X"DD",X"77",
		X"17",X"3A",X"05",X"4D",X"81",X"DD",X"77",X"16",X"3A",X"06",X"4D",X"2F",X"83",X"DD",X"77",X"19",
		X"3A",X"07",X"4D",X"81",X"DD",X"77",X"18",X"3A",X"08",X"4D",X"2F",X"83",X"DD",X"77",X"1B",X"3A",
		X"09",X"4D",X"81",X"DD",X"77",X"1A",X"3A",X"D2",X"4D",X"2F",X"83",X"DD",X"77",X"1D",X"3A",X"D3",
		X"4D",X"81",X"DD",X"77",X"1C",X"3A",X"A5",X"4D",X"A7",X"C2",X"94",X"17",X"3A",X"A4",X"4D",X"A7",
		X"C2",X"07",X"18",X"21",X"65",X"17",X"E5",X"3A",X"30",X"4D",X"E6",X"03",X"E7",X"E6",X"18",X"00",
		X"19",X"1A",X"19",X"38",X"19",X"F0",X"6A",X"F0",X"6A",X"F0",X"6A",X"F0",X"6A",X"F0",X"6A",X"F0",
		X"6A",X"F0",X"6A",X"F0",X"6A",X"78",X"A7",X"28",X"2B",X"0E",X"C0",X"3A",X"0A",X"4C",X"57",X"A1",
		X"20",X"05",X"7A",X"B1",X"C3",X"91",X"17",X"3A",X"30",X"4D",X"FE",X"02",X"20",X"09",X"CB",X"7A",
		X"28",X"12",X"7A",X"A9",X"C3",X"91",X"17",X"FE",X"03",X"20",X"09",X"CB",X"72",X"28",X"05",X"7A",
		X"A9",X"32",X"0A",X"4C",X"21",X"C0",X"4D",X"56",X"3E",X"1C",X"82",X"08",X"3A",X"70",X"4C",X"FE",
		X"03",X"CA",X"B1",X"17",X"08",X"DD",X"77",X"02",X"DD",X"77",X"04",X"DD",X"77",X"06",X"DD",X"77",
		X"08",X"0E",X"20",X"3A",X"AC",X"4D",X"A7",X"20",X"06",X"3A",X"A7",X"4D",X"A7",X"20",X"09",X"3A",
		X"2C",X"4D",X"87",X"82",X"81",X"DD",X"77",X"02",X"3A",X"AD",X"4D",X"A7",X"20",X"06",X"3A",X"A8",
		X"4D",X"A7",X"20",X"09",X"3A",X"2D",X"4D",X"87",X"82",X"81",X"DD",X"77",X"04",X"3A",X"AE",X"4D",
		X"A7",X"20",X"06",X"3A",X"A9",X"4D",X"A7",X"20",X"09",X"3A",X"2E",X"4D",X"87",X"82",X"81",X"DD",
		X"77",X"06",X"3A",X"AF",X"4D",X"A7",X"20",X"06",X"3A",X"AA",X"4D",X"A7",X"20",X"09",X"3A",X"2F",
		X"4D",X"87",X"82",X"81",X"DD",X"77",X"08",X"CD",X"3F",X"18",X"CD",X"87",X"18",X"CD",X"AC",X"18",
		X"78",X"A7",X"C8",X"0E",X"C0",X"3A",X"02",X"4C",X"B1",X"32",X"02",X"4C",X"3A",X"04",X"4C",X"B1",
		X"32",X"04",X"4C",X"3A",X"06",X"4C",X"B1",X"32",X"06",X"4C",X"3A",X"08",X"4C",X"B1",X"32",X"08",
		X"4C",X"3A",X"70",X"4C",X"FE",X"03",X"C8",X"3A",X"0C",X"4C",X"B1",X"32",X"0C",X"4C",X"C9",X"C9",
		X"3A",X"06",X"4E",X"D6",X"05",X"D8",X"3A",X"09",X"4D",X"E6",X"0F",X"FE",X"0C",X"38",X"04",X"16",
		X"18",X"18",X"12",X"FE",X"08",X"38",X"04",X"16",X"14",X"18",X"0A",X"FE",X"04",X"38",X"04",X"16",
		X"10",X"18",X"02",X"16",X"14",X"DD",X"72",X"04",X"14",X"DD",X"72",X"06",X"14",X"DD",X"72",X"08",
		X"14",X"DD",X"72",X"0C",X"DD",X"36",X"0A",X"3F",X"16",X"16",X"DD",X"72",X"05",X"DD",X"72",X"07",
		X"DD",X"72",X"09",X"DD",X"72",X"0D",X"C9",X"3A",X"07",X"4E",X"A7",X"C8",X"57",X"3A",X"3A",X"4D",
		X"D6",X"3D",X"20",X"04",X"DD",X"36",X"0B",X"00",X"7A",X"FE",X"0A",X"D8",X"DD",X"36",X"02",X"32",
		X"DD",X"36",X"03",X"1D",X"FE",X"0C",X"D8",X"DD",X"36",X"02",X"33",X"C9",X"3A",X"08",X"4E",X"A7",
		X"C8",X"57",X"3A",X"3A",X"4D",X"D6",X"3D",X"20",X"04",X"DD",X"36",X"0B",X"00",X"7A",X"FE",X"01",
		X"D8",X"3A",X"C0",X"4D",X"1E",X"08",X"83",X"DD",X"77",X"02",X"7A",X"FE",X"03",X"D8",X"3A",X"01",
		X"4D",X"E6",X"08",X"0F",X"0F",X"0F",X"1E",X"0A",X"83",X"DD",X"77",X"0C",X"3C",X"3C",X"DD",X"77",
		X"02",X"DD",X"36",X"0D",X"1F",X"C9",X"C3",X"1D",X"85",X"FE",X"04",X"38",X"05",X"DD",X"36",X"0A",
		X"2E",X"C9",X"FE",X"02",X"38",X"05",X"DD",X"36",X"0A",X"2C",X"C9",X"DD",X"36",X"0A",X"2E",X"C9",
		X"C3",X"32",X"85",X"FE",X"04",X"38",X"05",X"DD",X"36",X"0A",X"2D",X"C9",X"FE",X"02",X"38",X"05",
		X"DD",X"36",X"0A",X"2F",X"C9",X"DD",X"36",X"0A",X"30",X"C9",X"3A",X"09",X"4D",X"C3",X"46",X"85",
		X"1E",X"2E",X"CB",X"FB",X"DD",X"73",X"0A",X"C9",X"FE",X"04",X"38",X"04",X"1E",X"2C",X"18",X"F2",
		X"FE",X"02",X"30",X"EC",X"1E",X"30",X"18",X"EA",X"3A",X"08",X"4D",X"C3",X"5A",X"85",X"FE",X"04",
		X"38",X"08",X"1E",X"2F",X"CB",X"F3",X"DD",X"73",X"0A",X"C9",X"FE",X"02",X"38",X"44",X"1E",X"2D",
		X"18",X"F2",X"3A",X"70",X"4C",X"FE",X"02",X"28",X"08",X"FE",X"03",X"28",X"04",X"F1",X"F1",X"18",
		X"7B",X"F5",X"E5",X"D5",X"C5",X"21",X"64",X"80",X"22",X"08",X"4D",X"21",X"2C",X"2E",X"22",X"12",
		X"4D",X"22",X"39",X"4D",X"21",X"00",X"01",X"22",X"1C",X"4D",X"22",X"26",X"4D",X"3E",X"00",X"32",
		X"72",X"4C",X"3E",X"02",X"32",X"30",X"4D",X"32",X"3C",X"4D",X"CD",X"65",X"1D",X"C1",X"D1",X"E1",
		X"F1",X"C9",X"1E",X"2F",X"18",X"AE",X"06",X"04",X"ED",X"5B",X"39",X"4D",X"3A",X"AF",X"4D",X"A7",
		X"20",X"09",X"2A",X"37",X"4D",X"A7",X"ED",X"52",X"CA",X"DC",X"19",X"05",X"3A",X"AE",X"4D",X"A7",
		X"20",X"09",X"2A",X"35",X"4D",X"A7",X"ED",X"52",X"CA",X"DC",X"19",X"05",X"3A",X"AD",X"4D",X"A7",
		X"20",X"09",X"2A",X"33",X"4D",X"A7",X"ED",X"52",X"CA",X"DC",X"19",X"05",X"3A",X"AC",X"4D",X"A7",
		X"20",X"09",X"2A",X"31",X"4D",X"A7",X"ED",X"52",X"CC",X"52",X"19",X"05",X"78",X"32",X"A4",X"4D",
		X"32",X"A5",X"4D",X"A7",X"C8",X"21",X"A6",X"4D",X"5F",X"16",X"00",X"19",X"7E",X"A7",X"C8",X"AF",
		X"32",X"A5",X"4D",X"21",X"D0",X"4D",X"34",X"46",X"04",X"CD",X"90",X"28",X"21",X"BC",X"4E",X"CB",
		X"DE",X"C9",X"3A",X"A4",X"4D",X"A7",X"C0",X"3A",X"A6",X"4D",X"A7",X"C8",X"0E",X"04",X"06",X"04",
		X"DD",X"21",X"08",X"4D",X"3A",X"AF",X"4D",X"A7",X"20",X"13",X"3A",X"06",X"4D",X"DD",X"96",X"00",
		X"B9",X"30",X"0A",X"3A",X"07",X"4D",X"DD",X"96",X"01",X"B9",X"DA",X"DC",X"19",X"05",X"3A",X"AE",
		X"4D",X"A7",X"20",X"13",X"3A",X"04",X"4D",X"DD",X"96",X"00",X"B9",X"30",X"0A",X"3A",X"05",X"4D",
		X"DD",X"96",X"01",X"B9",X"DA",X"DC",X"19",X"05",X"3A",X"AD",X"4D",X"A7",X"20",X"13",X"3A",X"02",
		X"4D",X"DD",X"96",X"00",X"B9",X"30",X"0A",X"3A",X"03",X"4D",X"DD",X"96",X"01",X"B9",X"DA",X"DC",
		X"19",X"05",X"3A",X"AC",X"4D",X"A7",X"20",X"13",X"3A",X"00",X"4D",X"DD",X"96",X"00",X"B9",X"30",
		X"0A",X"3A",X"01",X"4D",X"DD",X"96",X"01",X"B9",X"DA",X"DC",X"19",X"05",X"C3",X"DC",X"19",X"3A",
		X"70",X"4C",X"FE",X"01",X"28",X"45",X"FE",X"02",X"28",X"41",X"FE",X"03",X"28",X"3D",X"21",X"9D",
		X"4D",X"3E",X"FF",X"BE",X"CA",X"99",X"1A",X"35",X"C9",X"3A",X"A6",X"4D",X"A7",X"CA",X"B7",X"1A",
		X"2A",X"4C",X"4D",X"29",X"22",X"4C",X"4D",X"2A",X"4A",X"4D",X"ED",X"6A",X"22",X"4A",X"4D",X"D0",
		X"21",X"4C",X"4D",X"34",X"C3",X"CB",X"1A",X"2A",X"48",X"4D",X"29",X"22",X"48",X"4D",X"2A",X"46",
		X"4D",X"ED",X"6A",X"22",X"46",X"4D",X"D0",X"21",X"48",X"4D",X"34",X"3A",X"0E",X"4E",X"32",X"9E",
		X"4D",X"3A",X"72",X"4E",X"4F",X"3A",X"09",X"4E",X"A1",X"4F",X"21",X"3A",X"4D",X"7E",X"06",X"21",
		X"90",X"38",X"09",X"7E",X"06",X"3B",X"90",X"30",X"03",X"C3",X"33",X"1B",X"3E",X"01",X"32",X"BF",
		X"4D",X"3A",X"00",X"4E",X"FE",X"01",X"CA",X"A8",X"1D",X"3A",X"04",X"4E",X"FE",X"10",X"D2",X"A8",
		X"1D",X"79",X"A7",X"28",X"06",X"3A",X"40",X"50",X"C3",X"0E",X"1B",X"3A",X"00",X"50",X"CB",X"4F",
		X"C2",X"21",X"1B",X"2A",X"89",X"32",X"3E",X"02",X"32",X"30",X"4D",X"22",X"1C",X"4D",X"C3",X"D8",
		X"1B",X"CB",X"57",X"C2",X"D8",X"1B",X"2A",X"85",X"32",X"AF",X"32",X"30",X"4D",X"22",X"1C",X"4D",
		X"C3",X"D8",X"1B",X"3A",X"00",X"4E",X"FE",X"01",X"CA",X"A8",X"1D",X"3A",X"04",X"4E",X"FE",X"10",
		X"D2",X"A8",X"1D",X"79",X"A7",X"28",X"06",X"3A",X"40",X"50",X"C3",X"50",X"1B",X"3A",X"00",X"50",
		X"CB",X"4F",X"CA",X"60",X"1E",X"CB",X"57",X"CA",X"70",X"1E",X"CB",X"47",X"CA",X"7F",X"1E",X"CB",
		X"5F",X"CA",X"8F",X"1E",X"2A",X"1C",X"4D",X"22",X"26",X"4D",X"06",X"01",X"DD",X"21",X"26",X"4D",
		X"FD",X"21",X"39",X"4D",X"CD",X"DC",X"1E",X"E6",X"C0",X"D6",X"C0",X"20",X"4B",X"05",X"C2",X"9E",
		X"1B",X"3A",X"30",X"4D",X"0F",X"DA",X"93",X"1B",X"3A",X"09",X"4D",X"E6",X"07",X"FE",X"04",X"C8",
		X"C3",X"C8",X"1B",X"3A",X"08",X"4D",X"E6",X"07",X"FE",X"04",X"C8",X"C3",X"C8",X"1B",X"DD",X"21",
		X"1C",X"4D",X"CD",X"DC",X"1E",X"E6",X"C0",X"D6",X"C0",X"20",X"2D",X"3A",X"30",X"4D",X"0F",X"DA",
		X"BD",X"1B",X"3A",X"09",X"4D",X"E6",X"07",X"FE",X"04",X"C8",X"C3",X"D8",X"1B",X"3A",X"08",X"4D",
		X"E6",X"07",X"FE",X"04",X"C8",X"C3",X"D8",X"1B",X"2A",X"26",X"4D",X"22",X"1C",X"4D",X"05",X"CA",
		X"D8",X"1B",X"3A",X"3C",X"4D",X"32",X"30",X"4D",X"DD",X"21",X"1C",X"4D",X"FD",X"21",X"08",X"4D",
		X"CD",X"CD",X"1E",X"3A",X"30",X"4D",X"0F",X"DA",X"FD",X"1B",X"7D",X"E6",X"07",X"FE",X"04",X"CA",
		X"0D",X"1C",X"DA",X"F9",X"1B",X"2D",X"C3",X"0D",X"1C",X"2C",X"C3",X"0D",X"1C",X"7C",X"E6",X"07",
		X"FE",X"04",X"CA",X"0D",X"1C",X"DA",X"0C",X"1C",X"25",X"C3",X"0D",X"1C",X"24",X"22",X"08",X"4D",
		X"CD",X"E5",X"1E",X"22",X"39",X"4D",X"DD",X"21",X"BF",X"4D",X"DD",X"7E",X"00",X"DD",X"36",X"00",
		X"00",X"A7",X"C0",X"3A",X"D2",X"4D",X"A7",X"28",X"29",X"3A",X"D4",X"4D",X"A7",X"28",X"23",X"08",
		X"3A",X"70",X"4C",X"FE",X"03",X"C8",X"08",X"2A",X"08",X"4D",X"11",X"94",X"80",X"C3",X"D3",X"86",
		X"06",X"19",X"4F",X"CD",X"42",X"00",X"CD",X"AF",X"11",X"F7",X"54",X"05",X"00",X"21",X"BC",X"4E",
		X"CB",X"D6",X"3E",X"FF",X"32",X"9D",X"4D",X"2A",X"39",X"4D",X"CD",X"69",X"00",X"7E",X"FE",X"10",
		X"28",X"43",X"FE",X"4D",X"CC",X"EE",X"1C",X"FE",X"14",X"CC",X"77",X"1D",X"28",X"37",X"FE",X"B0",
		X"D0",X"FE",X"90",X"D8",X"3A",X"FD",X"4D",X"3C",X"32",X"FD",X"4D",X"DD",X"21",X"00",X"4C",X"3E",
		X"1C",X"DD",X"BE",X"02",X"CA",X"90",X"B3",X"DD",X"BE",X"04",X"CA",X"90",X"B3",X"DD",X"BE",X"06",
		X"CA",X"90",X"B3",X"DD",X"BE",X"08",X"CA",X"90",X"B3",X"E5",X"CD",X"15",X"87",X"CD",X"90",X"B3",
		X"CD",X"69",X"B4",X"E1",X"C9",X"3A",X"72",X"4C",X"A7",X"28",X"08",X"3D",X"32",X"72",X"4C",X"A7",
		X"CC",X"65",X"1D",X"7E",X"DD",X"21",X"0E",X"4E",X"DD",X"34",X"00",X"E6",X"0F",X"CB",X"3F",X"06",
		X"40",X"70",X"06",X"19",X"4F",X"CB",X"39",X"CD",X"42",X"00",X"3C",X"FE",X"01",X"CA",X"D1",X"1C",
		X"87",X"32",X"9D",X"4D",X"CD",X"9F",X"1E",X"CD",X"F9",X"1D",X"21",X"BC",X"4E",X"3A",X"0E",X"4E",
		X"FE",X"04",X"DC",X"E3",X"B5",X"0F",X"DA",X"A3",X"1D",X"CB",X"C6",X"CB",X"8E",X"C9",X"F5",X"E5",
		X"3A",X"14",X"4E",X"A7",X"28",X"06",X"CD",X"65",X"1D",X"CD",X"5F",X"B6",X"E1",X"F1",X"C9",X"3A",
		X"13",X"4E",X"FE",X"01",X"D2",X"22",X"1D",X"3A",X"79",X"4C",X"FE",X"02",X"D2",X"22",X"1D",X"F5",
		X"EF",X"1C",X"36",X"EF",X"20",X"10",X"3A",X"79",X"4C",X"3C",X"32",X"79",X"4C",X"CD",X"30",X"05",
		X"F1",X"C9",X"3A",X"14",X"4E",X"FE",X"06",X"30",X"1D",X"3A",X"7A",X"4C",X"FE",X"02",X"D2",X"46",
		X"1D",X"3C",X"32",X"7A",X"4C",X"F5",X"EF",X"1C",X"36",X"EF",X"20",X"11",X"CD",X"00",X"87",X"21",
		X"9C",X"4E",X"CB",X"CE",X"F1",X"C9",X"F5",X"EF",X"1C",X"36",X"EF",X"20",X"12",X"21",X"BC",X"4E",
		X"CB",X"DE",X"F1",X"C9",X"F5",X"EF",X"1C",X"36",X"EF",X"20",X"13",X"EF",X"21",X"12",X"21",X"BC",
		X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"AF",X"32",X"72",X"4C",X"06",X"14",X"CD",
		X"DF",X"2A",X"E1",X"D1",X"C1",X"F1",X"C9",X"F5",X"E5",X"3A",X"70",X"4C",X"FE",X"03",X"28",X"07",
		X"3A",X"70",X"4C",X"FE",X"02",X"20",X"19",X"EF",X"1C",X"16",X"3E",X"02",X"32",X"CC",X"4E",X"32",
		X"DC",X"4E",X"3A",X"70",X"4C",X"FE",X"03",X"3E",X"20",X"20",X"02",X"3E",X"40",X"32",X"72",X"4C",
		X"E1",X"F1",X"C9",X"CB",X"86",X"CB",X"CE",X"C9",X"21",X"1C",X"4D",X"7E",X"A7",X"CA",X"BD",X"1D",
		X"3A",X"08",X"4D",X"E6",X"07",X"FE",X"04",X"CA",X"C7",X"1D",X"C3",X"EB",X"1D",X"3A",X"09",X"4D",
		X"E6",X"07",X"FE",X"04",X"C2",X"EB",X"1D",X"3E",X"05",X"CD",X"C8",X"A6",X"38",X"03",X"EF",X"17",
		X"00",X"DD",X"21",X"26",X"4D",X"FD",X"21",X"12",X"4D",X"CD",X"CD",X"1E",X"22",X"12",X"4D",X"2A",
		X"26",X"4D",X"22",X"1C",X"4D",X"3A",X"3C",X"4D",X"32",X"30",X"4D",X"DD",X"21",X"1C",X"4D",X"FD",
		X"21",X"08",X"4D",X"CD",X"CD",X"1E",X"C3",X"0D",X"1C",X"3A",X"9D",X"4D",X"FE",X"06",X"C0",X"2A",
		X"BD",X"4D",X"22",X"CB",X"4D",X"3E",X"01",X"32",X"A6",X"4D",X"32",X"A7",X"4D",X"32",X"A8",X"4D",
		X"32",X"A9",X"4D",X"32",X"AA",X"4D",X"32",X"B1",X"4D",X"32",X"B2",X"4D",X"32",X"B3",X"4D",X"32",
		X"B4",X"4D",X"32",X"B5",X"4D",X"AF",X"32",X"C8",X"4D",X"32",X"D0",X"4D",X"DD",X"21",X"00",X"4C",
		X"3A",X"70",X"4C",X"FE",X"03",X"CA",X"CE",X"B3",X"DD",X"36",X"02",X"1C",X"DD",X"36",X"04",X"1C",
		X"DD",X"36",X"06",X"1C",X"DD",X"36",X"08",X"1C",X"DD",X"36",X"03",X"11",X"DD",X"36",X"05",X"11",
		X"DD",X"36",X"07",X"11",X"DD",X"36",X"09",X"11",X"21",X"AC",X"4E",X"CB",X"EE",X"CB",X"BE",X"C9",
		X"2A",X"89",X"32",X"3E",X"02",X"32",X"3C",X"4D",X"22",X"26",X"4D",X"06",X"00",X"C3",X"6C",X"1B",
		X"2A",X"85",X"32",X"AF",X"32",X"3C",X"4D",X"22",X"26",X"4D",X"06",X"00",X"C3",X"6C",X"1B",X"2A",
		X"8B",X"32",X"3E",X"03",X"32",X"3C",X"4D",X"22",X"26",X"4D",X"06",X"00",X"C3",X"6C",X"1B",X"2A",
		X"87",X"32",X"3E",X"01",X"32",X"3C",X"4D",X"22",X"26",X"4D",X"06",X"00",X"C3",X"6C",X"1B",X"3A",
		X"12",X"4E",X"A7",X"CA",X"AB",X"1E",X"21",X"9F",X"4D",X"34",X"C9",X"3A",X"A3",X"4D",X"A7",X"C0",
		X"3A",X"A2",X"4D",X"A7",X"CA",X"BC",X"1E",X"21",X"11",X"4E",X"34",X"C9",X"3A",X"A1",X"4D",X"A7",
		X"CA",X"C8",X"1E",X"21",X"10",X"4E",X"34",X"C9",X"21",X"0F",X"4E",X"34",X"C9",X"FD",X"7E",X"00",
		X"DD",X"86",X"00",X"6F",X"FD",X"7E",X"01",X"DD",X"86",X"01",X"67",X"C9",X"CD",X"CD",X"1E",X"CD",
		X"69",X"00",X"7E",X"A7",X"C9",X"7D",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"20",X"6F",X"7C",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"1E",X"67",X"C9",X"F5",X"C5",X"7D",X"D6",X"20",X"6F",
		X"7C",X"D6",X"20",X"67",X"06",X"00",X"CB",X"24",X"CB",X"24",X"CB",X"24",X"CB",X"24",X"CB",X"10",
		X"CB",X"24",X"CB",X"10",X"4C",X"26",X"00",X"09",X"01",X"40",X"40",X"09",X"C1",X"F1",X"C9",X"CD",
		X"69",X"00",X"11",X"00",X"04",X"19",X"C9",X"CD",X"1F",X"1F",X"7E",X"FE",X"1B",X"C3",X"CE",X"35",
		X"AF",X"02",X"C9",X"3A",X"A1",X"4D",X"A7",X"C0",X"3A",X"12",X"4E",X"A7",X"CA",X"48",X"1F",X"3A",
		X"9F",X"4D",X"FE",X"07",X"C0",X"C3",X"50",X"1F",X"21",X"B8",X"4D",X"3A",X"0F",X"4E",X"BE",X"D8",
		X"3E",X"02",X"32",X"A1",X"4D",X"C9",X"3A",X"A2",X"4D",X"A7",X"C0",X"3A",X"12",X"4E",X"A7",X"CA",
		X"6B",X"1F",X"3A",X"9F",X"4D",X"FE",X"11",X"C0",X"C3",X"73",X"1F",X"21",X"B9",X"4D",X"3A",X"10",
		X"4E",X"BE",X"D8",X"3E",X"03",X"32",X"A2",X"4D",X"C9",X"3A",X"A3",X"4D",X"A7",X"C0",X"3A",X"12",
		X"4E",X"A7",X"CA",X"93",X"1F",X"3A",X"9F",X"4D",X"FE",X"20",X"C0",X"AF",X"32",X"12",X"4E",X"32",
		X"9F",X"4D",X"C9",X"21",X"BA",X"4D",X"3A",X"11",X"4E",X"BE",X"D8",X"3E",X"03",X"32",X"A3",X"4D",
		X"C9",X"3A",X"A3",X"4D",X"A7",X"C8",X"21",X"0E",X"4E",X"3A",X"B6",X"4D",X"A7",X"C2",X"BE",X"1F",
		X"3E",X"F4",X"96",X"47",X"3A",X"BB",X"4D",X"90",X"D8",X"3E",X"01",X"32",X"B6",X"4D",X"3A",X"B7",
		X"4D",X"A7",X"C0",X"3E",X"F4",X"96",X"47",X"3A",X"BC",X"4D",X"90",X"D8",X"3E",X"01",X"32",X"B7",
		X"4D",X"C9",X"20",X"96",X"01",X"ED",X"47",X"21",X"00",X"50",X"06",X"08",X"AF",X"77",X"2C",X"10",
		X"FC",X"21",X"00",X"60",X"7E",X"FE",X"4D",X"20",X"16",X"23",X"7E",X"FE",X"49",X"20",X"10",X"23",
		X"7E",X"FE",X"4B",X"20",X"0A",X"23",X"7E",X"FE",X"59",X"20",X"04",X"23",X"C3",X"7F",X"1A",X"AF",
		X"ED",X"47",X"21",X"00",X"50",X"06",X"08",X"AF",X"77",X"2C",X"10",X"FC",X"21",X"00",X"40",X"06",
		X"04",X"32",X"C0",X"50",X"32",X"07",X"50",X"3E",X"40",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F1",
		X"06",X"04",X"32",X"C0",X"50",X"AF",X"32",X"07",X"50",X"3E",X"0F",X"77",X"2C",X"20",X"FC",X"24",
		X"10",X"F0",X"ED",X"56",X"AF",X"32",X"07",X"50",X"3C",X"32",X"00",X"50",X"FB",X"76",X"C3",X"6C",
		X"00",X"21",X"04",X"4E",X"34",X"C9",X"78",X"E6",X"01",X"E7",X"4E",X"20",X"5B",X"20",X"3E",X"40",
		X"01",X"04",X"00",X"21",X"00",X"40",X"CF",X"0D",X"20",X"FC",X"C9",X"3E",X"40",X"21",X"40",X"40",
		X"01",X"04",X"80",X"CF",X"0D",X"20",X"FC",X"C9",X"AF",X"01",X"04",X"00",X"21",X"00",X"44",X"CF",
		X"0D",X"20",X"FC",X"C9",X"21",X"00",X"40",X"CD",X"0D",X"94",X"0A",X"A7",X"C8",X"FA",X"87",X"20",
		X"5F",X"16",X"00",X"19",X"2B",X"03",X"0A",X"23",X"77",X"F5",X"E5",X"11",X"E0",X"83",X"7D",X"E6",
		X"1F",X"87",X"26",X"00",X"6F",X"19",X"D1",X"A7",X"ED",X"52",X"F1",X"EE",X"01",X"77",X"EB",X"03",
		X"C3",X"7A",X"20",X"10",X"11",X"12",X"13",X"14",X"01",X"03",X"04",X"06",X"07",X"08",X"09",X"0A",
		X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"14",X"C0",X"50",X"80",X"50",X"C0",X"50",X"F5",X"08",
		X"F5",X"AF",X"32",X"00",X"50",X"F3",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"21",X"8C",X"4E",
		X"11",X"50",X"50",X"01",X"10",X"00",X"ED",X"B0",X"3A",X"CC",X"4E",X"A7",X"3A",X"CF",X"4E",X"20",
		X"03",X"3A",X"9F",X"4E",X"32",X"45",X"50",X"3A",X"DC",X"4E",X"A7",X"3A",X"DF",X"4E",X"20",X"03",
		X"3A",X"AF",X"4E",X"32",X"4A",X"50",X"3A",X"EC",X"4E",X"A7",X"3A",X"EF",X"4E",X"20",X"03",X"3A",
		X"BF",X"4E",X"32",X"4F",X"50",X"21",X"02",X"4C",X"11",X"22",X"4C",X"01",X"1C",X"00",X"ED",X"B0",
		X"DD",X"21",X"20",X"4C",X"DD",X"7E",X"02",X"07",X"07",X"DD",X"77",X"02",X"DD",X"7E",X"04",X"07",
		X"07",X"DD",X"77",X"04",X"DD",X"7E",X"06",X"07",X"07",X"DD",X"77",X"06",X"DD",X"7E",X"08",X"07",
		X"07",X"DD",X"77",X"08",X"DD",X"7E",X"0A",X"07",X"07",X"DD",X"77",X"0A",X"DD",X"7E",X"0C",X"07",
		X"07",X"DD",X"77",X"0C",X"3A",X"D1",X"4D",X"FE",X"01",X"20",X"38",X"DD",X"21",X"20",X"4C",X"3A",
		X"A4",X"4D",X"87",X"5F",X"16",X"00",X"DD",X"19",X"2A",X"24",X"4C",X"ED",X"5B",X"34",X"4C",X"DD",
		X"7E",X"00",X"32",X"24",X"4C",X"DD",X"7E",X"01",X"32",X"25",X"4C",X"DD",X"7E",X"10",X"32",X"34",
		X"4C",X"DD",X"7E",X"11",X"32",X"35",X"4C",X"DD",X"75",X"00",X"DD",X"74",X"01",X"DD",X"73",X"10",
		X"DD",X"72",X"11",X"3A",X"A6",X"4D",X"A7",X"CA",X"A6",X"21",X"ED",X"4B",X"22",X"4C",X"ED",X"5B",
		X"32",X"4C",X"2A",X"2A",X"4C",X"22",X"22",X"4C",X"2A",X"3A",X"4C",X"22",X"32",X"4C",X"ED",X"43",
		X"2A",X"4C",X"ED",X"53",X"3A",X"4C",X"21",X"22",X"4C",X"11",X"F2",X"4F",X"01",X"0E",X"00",X"ED",
		X"B0",X"21",X"32",X"4C",X"11",X"62",X"50",X"01",X"0E",X"00",X"ED",X"B0",X"3A",X"70",X"4C",X"FE",
		X"03",X"20",X"22",X"3A",X"FF",X"47",X"32",X"04",X"50",X"3C",X"E6",X"01",X"32",X"FF",X"47",X"32",
		X"05",X"50",X"E6",X"01",X"28",X"0F",X"3A",X"02",X"4E",X"A7",X"20",X"09",X"CD",X"B6",X"B0",X"CD",
		X"06",X"B1",X"CD",X"2D",X"B1",X"CD",X"10",X"04",X"CD",X"55",X"04",X"CD",X"30",X"06",X"3A",X"00",
		X"4E",X"A7",X"28",X"12",X"CD",X"04",X"06",X"CD",X"C7",X"16",X"CD",X"56",X"16",X"CD",X"B8",X"04",
		X"CD",X"FE",X"04",X"CD",X"64",X"05",X"3A",X"00",X"4E",X"3D",X"20",X"06",X"32",X"AC",X"4E",X"32",
		X"BC",X"4E",X"3E",X"55",X"47",X"CD",X"2C",X"AF",X"E6",X"0F",X"F6",X"FA",X"3C",X"C4",X"38",X"25",
		X"CD",X"B4",X"2B",X"CD",X"42",X"2B",X"3A",X"70",X"4C",X"FE",X"03",X"20",X"16",X"3A",X"FF",X"47",
		X"E6",X"01",X"28",X"0F",X"3A",X"02",X"4E",X"A7",X"20",X"09",X"CD",X"19",X"B1",X"CD",X"2D",X"B1",
		X"CD",X"DB",X"B0",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"3A",X"00",X"4E",X"A7",X"28",X"08",
		X"3A",X"40",X"50",X"E6",X"10",X"CA",X"00",X"00",X"3E",X"01",X"32",X"00",X"50",X"FB",X"F1",X"08",
		X"F1",X"C9",X"21",X"00",X"40",X"C3",X"3A",X"94",X"16",X"00",X"06",X"1E",X"0E",X"08",X"DD",X"7E",
		X"00",X"FD",X"5E",X"00",X"19",X"07",X"30",X"02",X"36",X"10",X"FD",X"23",X"0D",X"20",X"F2",X"DD",
		X"23",X"05",X"20",X"E8",X"21",X"34",X"4E",X"C3",X"D7",X"94",X"21",X"00",X"40",X"C3",X"3F",X"94",
		X"16",X"00",X"06",X"1E",X"0E",X"08",X"FD",X"5E",X"00",X"19",X"7E",X"FE",X"10",X"37",X"28",X"01",
		X"3F",X"DD",X"CB",X"00",X"16",X"FD",X"23",X"0D",X"20",X"EC",X"DD",X"23",X"05",X"20",X"E5",X"21",
		X"64",X"40",X"C3",X"05",X"95",X"21",X"16",X"4E",X"3E",X"FF",X"06",X"1E",X"CF",X"3E",X"14",X"06",
		X"04",X"CF",X"C9",X"58",X"78",X"FE",X"02",X"3E",X"1F",X"C3",X"99",X"95",X"10",X"21",X"40",X"44",
		X"01",X"04",X"80",X"CF",X"0D",X"20",X"FC",X"3E",X"0F",X"06",X"40",X"21",X"C0",X"47",X"CF",X"7B",
		X"FE",X"01",X"C0",X"3E",X"1A",X"C3",X"F1",X"95",X"06",X"06",X"DD",X"21",X"A0",X"45",X"DD",X"77",
		X"0C",X"DD",X"77",X"18",X"DD",X"19",X"10",X"F6",X"3E",X"1B",X"06",X"05",X"DD",X"21",X"40",X"44",
		X"DD",X"77",X"0E",X"DD",X"77",X"0F",X"DD",X"77",X"10",X"DD",X"19",X"10",X"F3",X"06",X"05",X"DD",
		X"21",X"20",X"47",X"DD",X"77",X"0E",X"DD",X"77",X"0F",X"DD",X"77",X"10",X"DD",X"19",X"10",X"F3",
		X"3E",X"18",X"32",X"ED",X"45",X"32",X"0D",X"46",X"C9",X"AF",X"32",X"04",X"50",X"32",X"05",X"50",
		X"32",X"FD",X"4D",X"DD",X"21",X"00",X"4C",X"DD",X"36",X"02",X"20",X"DD",X"36",X"04",X"20",X"DD",
		X"36",X"06",X"20",X"DD",X"36",X"08",X"20",X"DD",X"36",X"0A",X"2C",X"DD",X"36",X"03",X"01",X"DD",
		X"36",X"05",X"03",X"DD",X"36",X"07",X"05",X"DD",X"36",X"09",X"07",X"DD",X"36",X"0B",X"09",X"3A",
		X"70",X"4C",X"FE",X"03",X"20",X"0A",X"DD",X"36",X"0D",X"05",X"DD",X"36",X"0C",X"2C",X"18",X"08",
		X"DD",X"36",X"0D",X"09",X"DD",X"36",X"0C",X"0F",X"78",X"A7",X"C2",X"5E",X"24",X"21",X"64",X"80",
		X"22",X"00",X"4D",X"21",X"7C",X"80",X"22",X"02",X"4D",X"21",X"7C",X"90",X"22",X"04",X"4D",X"21",
		X"7C",X"70",X"22",X"06",X"4D",X"21",X"C4",X"70",X"22",X"08",X"4D",X"3A",X"70",X"4C",X"FE",X"03",
		X"28",X"06",X"21",X"C4",X"80",X"22",X"08",X"4D",X"21",X"2C",X"2E",X"22",X"0A",X"4D",X"22",X"31",
		X"4D",X"21",X"2F",X"2E",X"22",X"0C",X"4D",X"22",X"33",X"4D",X"21",X"2F",X"30",X"22",X"0E",X"4D",
		X"22",X"35",X"4D",X"21",X"2F",X"2C",X"22",X"10",X"4D",X"22",X"37",X"4D",X"21",X"38",X"2C",X"22",
		X"12",X"4D",X"22",X"39",X"4D",X"3A",X"70",X"4C",X"FE",X"03",X"28",X"12",X"21",X"38",X"2E",X"22",
		X"12",X"4D",X"22",X"39",X"4D",X"21",X"38",X"30",X"22",X"C6",X"4F",X"22",X"C8",X"4F",X"21",X"00",
		X"01",X"22",X"14",X"4D",X"22",X"1E",X"4D",X"21",X"01",X"00",X"22",X"16",X"4D",X"22",X"20",X"4D",
		X"21",X"FF",X"00",X"22",X"18",X"4D",X"22",X"22",X"4D",X"21",X"FF",X"00",X"22",X"1A",X"4D",X"22",
		X"24",X"4D",X"21",X"00",X"01",X"22",X"1C",X"4D",X"22",X"26",X"4D",X"21",X"00",X"FF",X"22",X"CA",
		X"4F",X"22",X"CC",X"4F",X"21",X"02",X"01",X"22",X"28",X"4D",X"22",X"2C",X"4D",X"21",X"03",X"03",
		X"22",X"2A",X"4D",X"22",X"2E",X"4D",X"3E",X"00",X"32",X"72",X"4C",X"3E",X"02",X"32",X"30",X"4D",
		X"32",X"3C",X"4D",X"3E",X"00",X"32",X"CE",X"4F",X"32",X"CF",X"4F",X"21",X"C4",X"90",X"22",X"D2",
		X"4D",X"3A",X"70",X"4C",X"FE",X"03",X"C8",X"21",X"00",X"00",X"22",X"D2",X"4D",X"C9",X"C9",X"21",
		X"00",X"00",X"22",X"D2",X"4D",X"22",X"08",X"4D",X"22",X"00",X"4D",X"22",X"02",X"4D",X"22",X"04",
		X"4D",X"22",X"06",X"4D",X"C9",X"3E",X"55",X"32",X"94",X"4D",X"05",X"C8",X"3E",X"01",X"32",X"A0",
		X"4D",X"C9",X"3E",X"01",X"32",X"00",X"4E",X"AF",X"32",X"01",X"4E",X"C9",X"AF",X"11",X"00",X"4D",
		X"21",X"00",X"4E",X"12",X"13",X"A7",X"ED",X"52",X"C2",X"90",X"24",X"C9",X"DD",X"21",X"36",X"41",
		X"3A",X"71",X"4E",X"E6",X"0F",X"C6",X"30",X"DD",X"77",X"00",X"3A",X"71",X"4E",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"C8",X"C6",X"30",X"DD",X"77",X"20",X"C9",X"DD",X"21",X"55",X"40",X"00",X"00",
		X"47",X"E6",X"0F",X"DD",X"77",X"00",X"78",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C8",X"DD",X"77",
		X"20",X"C9",X"3A",X"80",X"50",X"47",X"E6",X"03",X"C2",X"E0",X"24",X"21",X"6E",X"4E",X"36",X"FF",
		X"4F",X"1F",X"CE",X"00",X"32",X"6B",X"4E",X"E6",X"02",X"A9",X"32",X"6D",X"4E",X"78",X"0F",X"0F",
		X"E6",X"03",X"3C",X"FE",X"04",X"20",X"01",X"3C",X"32",X"6F",X"4E",X"78",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"03",X"21",X"34",X"25",X"D7",X"32",X"71",X"4E",X"78",X"07",X"2F",X"E6",X"01",X"32",X"75",
		X"4E",X"78",X"07",X"07",X"2F",X"E6",X"01",X"47",X"3A",X"70",X"4C",X"FE",X"03",X"21",X"4A",X"25",
		X"20",X"03",X"21",X"4E",X"25",X"DF",X"22",X"73",X"4E",X"3A",X"40",X"50",X"07",X"2F",X"E6",X"01",
		X"32",X"72",X"4E",X"C9",X"40",X"60",X"80",X"FF",X"2A",X"6A",X"4C",X"CB",X"BD",X"22",X"6A",X"4C",
		X"C9",X"2A",X"6A",X"4C",X"CB",X"FD",X"22",X"6A",X"4C",X"C9",X"66",X"01",X"66",X"01",X"93",X"01",
		X"93",X"01",X"3A",X"C1",X"4D",X"CB",X"47",X"C2",X"7A",X"25",X"3A",X"B6",X"4D",X"A7",X"20",X"1A",
		X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",X"2A",X"0A",X"4D",X"3A",X"2C",X"4D",X"CD",X"7A",X"95",
		X"CD",X"9C",X"27",X"22",X"1E",X"4D",X"32",X"2C",X"4D",X"C9",X"2A",X"0A",X"4D",X"ED",X"5B",X"39",
		X"4D",X"3A",X"2C",X"4D",X"CD",X"9C",X"27",X"22",X"1E",X"4D",X"32",X"2C",X"4D",X"C9",X"3A",X"C1",
		X"4D",X"CB",X"47",X"C2",X"B0",X"25",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",X"2A",X"0C",X"4D",
		X"3A",X"2D",X"4D",X"CD",X"7A",X"95",X"CD",X"9C",X"27",X"22",X"20",X"4D",X"32",X"2D",X"4D",X"C9",
		X"ED",X"5B",X"39",X"4D",X"2A",X"1C",X"4D",X"29",X"29",X"19",X"EB",X"2A",X"0C",X"4D",X"3A",X"2D",
		X"4D",X"CD",X"9C",X"27",X"22",X"20",X"4D",X"32",X"2D",X"4D",X"C9",X"3A",X"C1",X"4D",X"CB",X"47",
		X"C2",X"ED",X"25",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",X"2A",X"0E",X"4D",X"CD",X"72",X"95",
		X"11",X"40",X"20",X"CD",X"9C",X"27",X"22",X"22",X"4D",X"32",X"2E",X"4D",X"C9",X"ED",X"4B",X"0A",
		X"4D",X"ED",X"5B",X"39",X"4D",X"2A",X"1C",X"4D",X"29",X"19",X"7D",X"87",X"91",X"6F",X"7C",X"87",
		X"90",X"67",X"EB",X"2A",X"0E",X"4D",X"3A",X"2E",X"4D",X"CD",X"9C",X"27",X"22",X"22",X"4D",X"32",
		X"2E",X"4D",X"C9",X"3A",X"C1",X"4D",X"CB",X"47",X"C2",X"35",X"26",X"3A",X"04",X"4E",X"FE",X"03",
		X"20",X"13",X"2A",X"10",X"4D",X"CD",X"77",X"95",X"11",X"AE",X"3A",X"CD",X"9C",X"27",X"22",X"24",
		X"4D",X"32",X"2F",X"4D",X"C9",X"DD",X"21",X"39",X"4D",X"FD",X"21",X"10",X"4D",X"CD",X"20",X"28",
		X"11",X"40",X"00",X"A7",X"ED",X"52",X"DA",X"22",X"26",X"2A",X"10",X"4D",X"ED",X"5B",X"39",X"4D",
		X"3A",X"2F",X"4D",X"CD",X"9C",X"27",X"22",X"24",X"4D",X"32",X"2F",X"4D",X"C9",X"3A",X"AC",X"4D",
		X"A7",X"CA",X"77",X"26",X"11",X"2C",X"2E",X"2A",X"0A",X"4D",X"3A",X"2C",X"4D",X"CD",X"9C",X"27",
		X"22",X"1E",X"4D",X"32",X"2C",X"4D",X"C9",X"3E",X"01",X"32",X"DA",X"4F",X"2A",X"0A",X"4D",X"3A",
		X"2C",X"4D",X"CD",X"54",X"27",X"22",X"1E",X"4D",X"32",X"2C",X"4D",X"C9",X"3A",X"AD",X"4D",X"A7",
		X"CA",X"A6",X"26",X"11",X"2C",X"2E",X"2A",X"0C",X"4D",X"3A",X"2D",X"4D",X"CD",X"9C",X"27",X"22",
		X"20",X"4D",X"32",X"2D",X"4D",X"C9",X"3E",X"02",X"32",X"DA",X"4F",X"2A",X"0C",X"4D",X"3A",X"2D",
		X"4D",X"CD",X"54",X"27",X"22",X"20",X"4D",X"32",X"2D",X"4D",X"C9",X"3A",X"AE",X"4D",X"A7",X"CA",
		X"D5",X"26",X"11",X"2C",X"2E",X"2A",X"0E",X"4D",X"3A",X"2E",X"4D",X"CD",X"9C",X"27",X"22",X"22",
		X"4D",X"32",X"2E",X"4D",X"C9",X"3E",X"03",X"32",X"DA",X"4F",X"2A",X"0E",X"4D",X"3A",X"2E",X"4D",
		X"CD",X"54",X"27",X"22",X"22",X"4D",X"32",X"2E",X"4D",X"C9",X"3A",X"AF",X"4D",X"A7",X"CA",X"04",
		X"27",X"11",X"2C",X"2E",X"2A",X"10",X"4D",X"3A",X"2F",X"4D",X"CD",X"9C",X"27",X"22",X"24",X"4D",
		X"32",X"2F",X"4D",X"C9",X"3E",X"04",X"32",X"DA",X"4F",X"2A",X"10",X"4D",X"3A",X"2F",X"4D",X"CD",
		X"54",X"27",X"22",X"24",X"4D",X"32",X"2F",X"4D",X"C9",X"3A",X"A7",X"4D",X"A7",X"CA",X"34",X"27",
		X"2A",X"12",X"4D",X"ED",X"5B",X"0C",X"4D",X"3A",X"3C",X"4D",X"CD",X"9C",X"27",X"22",X"26",X"4D",
		X"32",X"3C",X"4D",X"C9",X"2A",X"39",X"4D",X"ED",X"4B",X"0C",X"4D",X"7D",X"87",X"91",X"6F",X"7C",
		X"87",X"90",X"67",X"EB",X"2A",X"12",X"4D",X"3A",X"3C",X"4D",X"CD",X"9C",X"27",X"22",X"26",X"4D",
		X"32",X"3C",X"4D",X"C9",X"22",X"3E",X"4D",X"EE",X"02",X"32",X"3D",X"4D",X"CD",X"59",X"28",X"E6",
		X"03",X"21",X"3B",X"4D",X"77",X"87",X"5F",X"16",X"00",X"DD",X"21",X"85",X"32",X"DD",X"19",X"FD",
		X"21",X"3E",X"4D",X"3A",X"3D",X"4D",X"BE",X"CA",X"8D",X"27",X"CD",X"DC",X"1E",X"E6",X"C0",X"D6",
		X"C0",X"28",X"0A",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"3A",X"3B",X"4D",X"C9",X"DD",X"23",X"DD",
		X"23",X"21",X"3B",X"4D",X"7E",X"3C",X"E6",X"03",X"77",X"C3",X"73",X"27",X"22",X"3E",X"4D",X"ED",
		X"53",X"40",X"4D",X"32",X"3B",X"4D",X"EE",X"02",X"32",X"3D",X"4D",X"21",X"FF",X"FF",X"22",X"44",
		X"4D",X"DD",X"21",X"85",X"32",X"FD",X"21",X"3E",X"4D",X"21",X"C7",X"4D",X"36",X"00",X"3A",X"3D",
		X"4D",X"BE",X"CA",X"FC",X"27",X"CD",X"CD",X"1E",X"22",X"42",X"4D",X"CD",X"69",X"00",X"7E",X"E6",
		X"C0",X"D6",X"C0",X"28",X"27",X"DD",X"E5",X"FD",X"E5",X"DD",X"21",X"40",X"4D",X"FD",X"21",X"42",
		X"4D",X"CD",X"20",X"28",X"FD",X"E1",X"DD",X"E1",X"EB",X"2A",X"44",X"4D",X"A7",X"ED",X"52",X"DA",
		X"FC",X"27",X"ED",X"53",X"44",X"4D",X"3A",X"C7",X"4D",X"32",X"3B",X"4D",X"DD",X"23",X"DD",X"23",
		X"21",X"C7",X"4D",X"34",X"3E",X"04",X"BE",X"C2",X"BE",X"27",X"3A",X"3B",X"4D",X"87",X"5F",X"16",
		X"00",X"DD",X"21",X"85",X"32",X"DD",X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"CB",X"3F",X"C9",
		X"DD",X"7E",X"00",X"FD",X"46",X"00",X"90",X"D2",X"2F",X"28",X"78",X"DD",X"46",X"00",X"90",X"CD",
		X"48",X"28",X"E5",X"DD",X"7E",X"01",X"FD",X"46",X"01",X"90",X"D2",X"42",X"28",X"78",X"DD",X"46",
		X"01",X"90",X"CD",X"48",X"28",X"C1",X"09",X"C9",X"67",X"5F",X"2E",X"00",X"55",X"0E",X"08",X"29",
		X"D2",X"54",X"28",X"19",X"0D",X"C2",X"4F",X"28",X"C9",X"2A",X"C9",X"4D",X"54",X"5D",X"29",X"29",
		X"19",X"23",X"7C",X"E6",X"1F",X"67",X"7E",X"22",X"C9",X"4D",X"C9",X"11",X"40",X"40",X"21",X"C0",
		X"43",X"A7",X"ED",X"52",X"C8",X"1A",X"FE",X"10",X"CA",X"89",X"28",X"FE",X"12",X"CA",X"89",X"28",
		X"FE",X"14",X"CA",X"89",X"28",X"13",X"C3",X"6E",X"28",X"3E",X"40",X"12",X"13",X"C3",X"6E",X"28",
		X"3A",X"00",X"4E",X"FE",X"01",X"C8",X"21",X"70",X"29",X"DF",X"EB",X"CD",X"64",X"29",X"7B",X"86",
		X"27",X"77",X"23",X"7A",X"8E",X"27",X"77",X"5F",X"23",X"3E",X"00",X"8E",X"27",X"77",X"57",X"EB",
		X"29",X"29",X"29",X"29",X"3A",X"71",X"4E",X"3D",X"BC",X"DC",X"AA",X"29",X"CD",X"EC",X"28",X"13",
		X"13",X"13",X"21",X"8A",X"4E",X"06",X"03",X"1A",X"BE",X"D8",X"20",X"05",X"1B",X"2B",X"10",X"F7",
		X"C9",X"3A",X"09",X"4E",X"3C",X"32",X"FE",X"4D",X"CD",X"64",X"29",X"11",X"88",X"4E",X"01",X"03",
		X"00",X"ED",X"B0",X"1B",X"01",X"04",X"03",X"21",X"F2",X"43",X"18",X"0F",X"3A",X"09",X"4E",X"01",
		X"04",X"03",X"21",X"FC",X"43",X"A7",X"28",X"03",X"21",X"E9",X"43",X"1A",X"0F",X"0F",X"0F",X"0F",
		X"CD",X"0B",X"29",X"1A",X"CD",X"0B",X"29",X"1B",X"10",X"F1",X"C9",X"E6",X"0F",X"28",X"04",X"0E",
		X"00",X"18",X"07",X"79",X"A7",X"28",X"03",X"3E",X"40",X"0D",X"77",X"2B",X"C9",X"21",X"E8",X"4D",
		X"23",X"23",X"7E",X"FE",X"4D",X"20",X"17",X"23",X"7E",X"FE",X"49",X"20",X"11",X"23",X"7E",X"FE",
		X"4B",X"20",X"0B",X"23",X"7E",X"FE",X"59",X"20",X"05",X"06",X"00",X"CD",X"DF",X"2A",X"AF",X"21",
		X"80",X"4E",X"06",X"08",X"CF",X"01",X"04",X"03",X"11",X"82",X"4E",X"21",X"FC",X"43",X"CD",X"FB",
		X"28",X"01",X"04",X"03",X"11",X"86",X"4E",X"21",X"E9",X"43",X"3A",X"70",X"4E",X"A7",X"20",X"9B",
		X"0E",X"06",X"18",X"97",X"3A",X"09",X"4E",X"21",X"80",X"4E",X"A7",X"C8",X"21",X"84",X"4E",X"C9",
		X"10",X"00",X"50",X"00",X"00",X"02",X"00",X"04",X"00",X"08",X"00",X"16",X"00",X"01",X"00",X"02",
		X"00",X"05",X"00",X"07",X"00",X"10",X"00",X"42",X"70",X"29",X"00",X"44",X"70",X"29",X"00",X"44",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"07",
		X"00",X"08",X"00",X"50",X"00",X"20",X"00",X"50",X"00",X"50",X"13",X"6B",X"62",X"1B",X"CB",X"46",
		X"C0",X"CB",X"C6",X"3E",X"01",X"32",X"CC",X"4E",X"32",X"DC",X"4E",X"21",X"14",X"4E",X"34",X"21",
		X"15",X"4E",X"34",X"46",X"21",X"1A",X"40",X"0E",X"05",X"78",X"A7",X"28",X"0E",X"FE",X"06",X"30",
		X"0A",X"3E",X"20",X"CD",X"09",X"2A",X"2B",X"2B",X"0D",X"10",X"F6",X"0D",X"F8",X"CD",X"F8",X"29",
		X"2B",X"2B",X"18",X"F7",X"3A",X"00",X"4E",X"FE",X"01",X"C8",X"CD",X"47",X"2A",X"12",X"44",X"09",
		X"0A",X"02",X"21",X"15",X"4E",X"46",X"18",X"CC",X"3E",X"40",X"E5",X"D5",X"77",X"23",X"77",X"11",
		X"1F",X"00",X"19",X"77",X"23",X"77",X"D1",X"E1",X"C9",X"E5",X"D5",X"11",X"1F",X"00",X"77",X"3C",
		X"23",X"77",X"3C",X"19",X"77",X"3C",X"23",X"77",X"D1",X"E1",X"C9",X"3A",X"6E",X"4E",X"FE",X"FF",
		X"20",X"05",X"06",X"02",X"C3",X"DF",X"2A",X"06",X"01",X"CD",X"DF",X"2A",X"3A",X"6E",X"4E",X"E6",
		X"F0",X"28",X"09",X"0F",X"0F",X"0F",X"0F",X"C6",X"30",X"32",X"34",X"40",X"3A",X"6E",X"4E",X"E6",
		X"0F",X"C6",X"30",X"32",X"33",X"40",X"C9",X"E1",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"23",
		X"7E",X"23",X"E5",X"EB",X"11",X"20",X"00",X"E5",X"C5",X"71",X"23",X"10",X"FC",X"C1",X"E1",X"19",
		X"3D",X"20",X"F4",X"C9",X"3A",X"00",X"4E",X"FE",X"01",X"C8",X"3A",X"13",X"4E",X"3C",X"FE",X"08",
		X"DA",X"75",X"2A",X"3E",X"07",X"11",X"76",X"3A",X"47",X"0E",X"07",X"21",X"04",X"40",X"1A",X"CD",
		X"09",X"2A",X"3E",X"04",X"84",X"67",X"13",X"1A",X"CD",X"FA",X"29",X"3E",X"FC",X"84",X"67",X"13",
		X"23",X"23",X"0D",X"10",X"E9",X"0D",X"F8",X"CD",X"F8",X"29",X"3E",X"04",X"84",X"67",X"AF",X"CD",
		X"FA",X"29",X"3E",X"FC",X"84",X"67",X"23",X"23",X"18",X"EB",X"FE",X"13",X"38",X"02",X"3E",X"13",
		X"D6",X"07",X"4F",X"06",X"00",X"21",X"76",X"3A",X"09",X"09",X"EB",X"06",X"07",X"C3",X"79",X"2A",
		X"47",X"E6",X"0F",X"C6",X"00",X"27",X"4F",X"78",X"E6",X"F0",X"28",X"0B",X"0F",X"0F",X"0F",X"0F",
		X"47",X"AF",X"C6",X"16",X"27",X"10",X"FB",X"81",X"27",X"C9",X"21",X"84",X"39",X"18",X"03",X"21",
		X"04",X"36",X"DF",X"5E",X"23",X"56",X"DD",X"21",X"00",X"44",X"DD",X"19",X"DD",X"E5",X"11",X"00",
		X"FC",X"DD",X"19",X"11",X"FF",X"FF",X"CB",X"7E",X"20",X"03",X"11",X"E0",X"FF",X"23",X"78",X"01",
		X"00",X"00",X"87",X"38",X"28",X"7E",X"FE",X"2F",X"28",X"09",X"DD",X"77",X"00",X"23",X"DD",X"19",
		X"04",X"18",X"F2",X"23",X"DD",X"E1",X"7E",X"A7",X"FA",X"25",X"2B",X"7E",X"DD",X"77",X"00",X"23",
		X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"77",X"00",X"DD",X"19",X"10",X"F9",X"C9",X"7E",X"FE",X"2F",
		X"28",X"0A",X"DD",X"36",X"00",X"40",X"23",X"DD",X"19",X"04",X"18",X"F1",X"23",X"04",X"ED",X"B1",
		X"18",X"D2",X"3A",X"00",X"4F",X"FE",X"00",X"28",X"0B",X"11",X"02",X"4C",X"21",X"50",X"4F",X"01",
		X"0E",X"00",X"ED",X"B0",X"3A",X"09",X"4E",X"21",X"72",X"4E",X"A6",X"28",X"0C",X"3A",X"0A",X"4C",
		X"FE",X"3F",X"20",X"05",X"3E",X"FF",X"32",X"0A",X"4C",X"21",X"26",X"A7",X"DD",X"21",X"CC",X"4E",
		X"FD",X"21",X"8C",X"4E",X"CD",X"EC",X"2B",X"47",X"3A",X"CC",X"4E",X"A7",X"28",X"04",X"78",X"32",
		X"91",X"4E",X"21",X"F6",X"A6",X"DD",X"21",X"DC",X"4E",X"FD",X"21",X"92",X"4E",X"CD",X"EC",X"2B",
		X"47",X"3A",X"DC",X"4E",X"A7",X"28",X"04",X"78",X"32",X"96",X"4E",X"21",X"5A",X"A7",X"DD",X"21",
		X"EC",X"4E",X"FD",X"21",X"97",X"4E",X"CD",X"EC",X"2B",X"47",X"3A",X"EC",X"4E",X"A7",X"C8",X"78",
		X"32",X"9B",X"4E",X"C9",X"21",X"9E",X"3A",X"DD",X"21",X"9C",X"4E",X"FD",X"21",X"8C",X"4E",X"CD",
		X"B1",X"2C",X"32",X"91",X"4E",X"21",X"AE",X"3A",X"DD",X"21",X"AC",X"4E",X"FD",X"21",X"92",X"4E",
		X"CD",X"B1",X"2C",X"32",X"96",X"4E",X"21",X"EE",X"3A",X"DD",X"21",X"BC",X"4E",X"FD",X"21",X"97",
		X"4E",X"CD",X"B1",X"2C",X"32",X"9B",X"4E",X"AF",X"32",X"90",X"4E",X"C9",X"DD",X"7E",X"00",X"A7",
		X"CA",X"B7",X"2C",X"4F",X"06",X"08",X"1E",X"80",X"7B",X"A1",X"20",X"05",X"CB",X"3B",X"10",X"F8",
		X"C9",X"DD",X"7E",X"02",X"A3",X"20",X"06",X"DD",X"73",X"02",X"C3",X"B8",X"35",X"DD",X"35",X"0C",
		X"C2",X"9A",X"2C",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",
		X"07",X"FE",X"F0",X"38",X"27",X"21",X"13",X"2C",X"E5",X"E6",X"0F",X"E7",X"18",X"2E",X"28",X"2E",
		X"3A",X"2E",X"4C",X"2E",X"5E",X"2E",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
		X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"70",X"2E",X"47",X"E6",X"1F",X"28",
		X"03",X"DD",X"70",X"0D",X"DD",X"4E",X"09",X"DD",X"7E",X"0B",X"E6",X"08",X"28",X"02",X"0E",X"00",
		X"DD",X"71",X"0F",X"78",X"07",X"07",X"07",X"E6",X"07",X"21",X"1E",X"3B",X"D7",X"DD",X"77",X"0C",
		X"08",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"FE",X"F5",X"20",X"10",X"23",X"DD",X"75",X"06",
		X"DD",X"74",X"07",X"08",X"CB",X"3F",X"DD",X"86",X"0C",X"DD",X"77",X"0C",X"78",X"E6",X"1F",X"28",
		X"09",X"E6",X"0F",X"21",X"2D",X"3B",X"D7",X"DD",X"77",X"0E",X"DD",X"6E",X"0E",X"26",X"00",X"DD",
		X"7E",X"0D",X"E6",X"10",X"28",X"02",X"3E",X"01",X"DD",X"86",X"04",X"CA",X"AB",X"2D",X"C3",X"A7",
		X"2D",X"DD",X"7E",X"00",X"A7",X"20",X"27",X"DD",X"7E",X"02",X"A7",X"C8",X"DD",X"36",X"02",X"00",
		X"DD",X"36",X"0D",X"00",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"00",X"FD",X"36",X"00",X"00",
		X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"00",X"FD",X"36",X"03",X"00",X"AF",X"C9",X"4F",X"06",
		X"08",X"1E",X"80",X"7B",X"A1",X"20",X"05",X"CB",X"3B",X"10",X"F8",X"C9",X"DD",X"7E",X"02",X"A3",
		X"20",X"3F",X"DD",X"73",X"02",X"05",X"78",X"07",X"07",X"07",X"4F",X"06",X"00",X"E5",X"09",X"DD",
		X"E5",X"D1",X"13",X"13",X"13",X"01",X"08",X"00",X"ED",X"B0",X"E1",X"DD",X"7E",X"06",X"E6",X"7F",
		X"DD",X"77",X"0C",X"DD",X"7E",X"04",X"DD",X"77",X"0E",X"DD",X"7E",X"09",X"47",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"DD",X"77",X"0B",X"E6",X"08",X"20",X"07",X"DD",X"70",X"0F",X"DD",X"36",X"0D",
		X"00",X"DD",X"35",X"0C",X"20",X"5A",X"DD",X"7E",X"08",X"A7",X"28",X"10",X"DD",X"35",X"08",X"20",
		X"0B",X"7B",X"2F",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C3",X"B1",X"2C",X"DD",X"7E",X"06",X"E6",
		X"7F",X"DD",X"77",X"0C",X"DD",X"CB",X"06",X"7E",X"28",X"16",X"DD",X"7E",X"05",X"ED",X"44",X"DD",
		X"77",X"05",X"DD",X"CB",X"0D",X"46",X"DD",X"CB",X"0D",X"C6",X"28",X"24",X"DD",X"CB",X"0D",X"86",
		X"DD",X"7E",X"04",X"DD",X"86",X"07",X"DD",X"77",X"04",X"DD",X"77",X"0E",X"DD",X"7E",X"09",X"DD",
		X"86",X"0A",X"DD",X"77",X"09",X"47",X"DD",X"7E",X"0B",X"E6",X"08",X"20",X"03",X"DD",X"70",X"0F",
		X"DD",X"7E",X"0E",X"DD",X"86",X"05",X"DD",X"77",X"0E",X"6F",X"26",X"00",X"DD",X"7E",X"03",X"E6",
		X"70",X"28",X"08",X"0F",X"0F",X"0F",X"0F",X"47",X"29",X"10",X"FD",X"FD",X"75",X"00",X"7D",X"0F",
		X"0F",X"0F",X"0F",X"FD",X"77",X"01",X"FD",X"74",X"02",X"7C",X"0F",X"0F",X"0F",X"0F",X"FD",X"77",
		X"03",X"DD",X"7E",X"0B",X"E7",X"E5",X"2D",X"E9",X"2D",X"EE",X"2D",X"FF",X"2D",X"06",X"2E",X"0D",
		X"2E",X"0E",X"2E",X"0F",X"2E",X"10",X"2E",X"11",X"2E",X"12",X"2E",X"13",X"2E",X"14",X"2E",X"15",
		X"2E",X"16",X"2E",X"17",X"2E",X"DD",X"7E",X"0F",X"C9",X"DD",X"7E",X"0F",X"18",X"09",X"3A",X"84",
		X"4C",X"E6",X"01",X"DD",X"7E",X"0F",X"C0",X"E6",X"0F",X"C8",X"3D",X"DD",X"77",X"0F",X"C9",X"3A",
		X"84",X"4C",X"E6",X"03",X"18",X"ED",X"3A",X"84",X"4C",X"E6",X"07",X"18",X"E6",X"C9",X"C9",X"C9",
		X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"DD",
		X"77",X"06",X"23",X"7E",X"DD",X"77",X"07",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"23",
		X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"03",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",
		X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"04",X"C9",X"DD",X"6E",X"06",X"DD",
		X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"09",X"C9",X"DD",X"6E",
		X"06",X"DD",X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"0B",X"C9",
		X"DD",X"7E",X"02",X"2F",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C3",X"B7",X"2C",X"3A",X"B1",X"4D",
		X"A7",X"C8",X"AF",X"32",X"B1",X"4D",X"21",X"85",X"32",X"3A",X"28",X"4D",X"EE",X"02",X"32",X"2C",
		X"4D",X"47",X"DF",X"22",X"1E",X"4D",X"3A",X"02",X"4E",X"FE",X"27",X"C0",X"22",X"14",X"4D",X"78",
		X"32",X"28",X"4D",X"C9",X"3A",X"B2",X"4D",X"A7",X"C8",X"AF",X"32",X"B2",X"4D",X"21",X"85",X"32",
		X"3A",X"29",X"4D",X"EE",X"02",X"32",X"2D",X"4D",X"47",X"DF",X"22",X"20",X"4D",X"3A",X"02",X"4E",
		X"FE",X"27",X"C0",X"22",X"16",X"4D",X"78",X"32",X"29",X"4D",X"C9",X"3A",X"B3",X"4D",X"A7",X"C8",
		X"AF",X"32",X"B3",X"4D",X"21",X"85",X"32",X"3A",X"2A",X"4D",X"EE",X"02",X"32",X"2E",X"4D",X"47",
		X"DF",X"22",X"22",X"4D",X"3A",X"02",X"4E",X"FE",X"27",X"C0",X"22",X"18",X"4D",X"78",X"32",X"2A",
		X"4D",X"C9",X"3A",X"B4",X"4D",X"A7",X"C8",X"AF",X"32",X"B4",X"4D",X"21",X"85",X"32",X"3A",X"2B",
		X"4D",X"EE",X"02",X"32",X"2F",X"4D",X"47",X"DF",X"22",X"24",X"4D",X"3A",X"02",X"4E",X"FE",X"27",
		X"C0",X"22",X"1A",X"4D",X"78",X"32",X"2B",X"4D",X"C9",X"F5",X"08",X"F5",X"ED",X"57",X"B7",X"28",
		X"06",X"F1",X"08",X"F1",X"C3",X"BE",X"20",X"F1",X"08",X"F1",X"C3",X"2D",X"2F",X"21",X"00",X"00",
		X"01",X"00",X"10",X"32",X"C0",X"50",X"79",X"86",X"4F",X"7D",X"C6",X"02",X"6F",X"FE",X"02",X"D2",
		X"36",X"2F",X"24",X"10",X"EE",X"79",X"A7",X"32",X"07",X"50",X"7C",X"FE",X"30",X"C2",X"30",X"2F",
		X"26",X"00",X"2C",X"7D",X"FE",X"02",X"DA",X"30",X"2F",X"C3",X"6D",X"2F",X"25",X"7C",X"E6",X"F0",
		X"32",X"07",X"50",X"0F",X"0F",X"0F",X"0F",X"5F",X"06",X"00",X"C3",X"E8",X"2F",X"31",X"9B",X"30",
		X"06",X"FF",X"E1",X"D1",X"48",X"32",X"C0",X"50",X"79",X"A3",X"77",X"C6",X"33",X"4F",X"2C",X"7D",
		X"E6",X"0F",X"C2",X"78",X"2F",X"79",X"87",X"87",X"81",X"C6",X"31",X"4F",X"7D",X"A7",X"C2",X"78",
		X"2F",X"24",X"15",X"C2",X"75",X"2F",X"3B",X"3B",X"3B",X"3B",X"E1",X"D1",X"48",X"32",X"C0",X"50",
		X"79",X"A3",X"4F",X"7E",X"A3",X"B9",X"C2",X"E0",X"2F",X"C6",X"33",X"4F",X"2C",X"7D",X"E6",X"0F",
		X"C2",X"A0",X"2F",X"79",X"87",X"87",X"81",X"C6",X"31",X"4F",X"7D",X"A7",X"C2",X"A0",X"2F",X"24",
		X"15",X"C2",X"9D",X"2F",X"3B",X"3B",X"3B",X"3B",X"78",X"D6",X"10",X"47",X"10",X"A4",X"F1",X"D1",
		X"FE",X"44",X"C2",X"70",X"2F",X"7B",X"EE",X"F0",X"C2",X"70",X"2F",X"06",X"01",X"C3",X"E8",X"2F",
		X"7B",X"E6",X"01",X"EE",X"01",X"5F",X"06",X"00",X"31",X"C0",X"4F",X"D9",X"21",X"00",X"4C",X"06",
		X"04",X"32",X"C0",X"50",X"36",X"00",X"2C",X"20",X"FB",X"24",X"10",X"F5",X"21",X"00",X"40",X"06",
		X"04",X"32",X"C0",X"50",X"3E",X"40",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F4",X"06",X"04",X"32",
		X"C0",X"50",X"3E",X"0F",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F4",X"D9",X"10",X"24",X"3E",X"0F",
		X"11",X"02",X"18",X"CD",X"AB",X"01",X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",X"41",X"40",X"56",
		X"4F",X"4C",X"41",X"54",X"49",X"4C",X"40",X"4F",X"4B",X"00",X"06",X"23",X"CD",X"DF",X"2A",X"C3",
		X"BB",X"30",X"7B",X"C6",X"30",X"32",X"84",X"41",X"C5",X"E5",X"06",X"24",X"CD",X"DF",X"2A",X"E1",
		X"7C",X"FE",X"40",X"2A",X"B3",X"30",X"38",X"11",X"FE",X"4C",X"2A",X"B5",X"30",X"30",X"0A",X"FE",
		X"44",X"2A",X"B7",X"30",X"38",X"03",X"2A",X"B9",X"30",X"7D",X"32",X"04",X"42",X"7C",X"32",X"64",
		X"42",X"3A",X"00",X"50",X"47",X"3A",X"40",X"50",X"B0",X"E6",X"01",X"20",X"11",X"C1",X"79",X"E6",
		X"0F",X"47",X"79",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"4F",X"ED",X"43",X"85",X"41",X"32",X"C0",
		X"50",X"3A",X"80",X"50",X"E6",X"08",X"28",X"F6",X"C3",X"D5",X"1F",X"00",X"4C",X"0F",X"04",X"00",
		X"4C",X"F0",X"04",X"00",X"40",X"0F",X"04",X"00",X"40",X"F0",X"04",X"00",X"44",X"0F",X"04",X"00",
		X"44",X"F0",X"04",X"4F",X"40",X"41",X"57",X"41",X"56",X"41",X"43",X"21",X"06",X"50",X"3E",X"01",
		X"77",X"2D",X"20",X"FC",X"AF",X"32",X"03",X"50",X"D6",X"04",X"ED",X"47",X"31",X"C0",X"4F",X"32",
		X"C0",X"50",X"AF",X"32",X"00",X"4E",X"3C",X"32",X"01",X"4E",X"32",X"00",X"50",X"FB",X"3A",X"00",
		X"50",X"2F",X"47",X"E6",X"A7",X"28",X"05",X"3E",X"02",X"32",X"9C",X"4E",X"3A",X"40",X"50",X"2F",
		X"4F",X"E6",X"27",X"28",X"05",X"3E",X"01",X"32",X"9C",X"4E",X"78",X"B1",X"E6",X"01",X"28",X"05",
		X"3E",X"08",X"32",X"BC",X"4E",X"78",X"B1",X"E6",X"02",X"28",X"05",X"3E",X"04",X"32",X"BC",X"4E",
		X"78",X"B1",X"E6",X"04",X"28",X"05",X"3E",X"10",X"32",X"BC",X"4E",X"78",X"B1",X"E6",X"08",X"28",
		X"05",X"3E",X"20",X"32",X"BC",X"4E",X"3A",X"80",X"50",X"E6",X"03",X"C6",X"25",X"47",X"CD",X"DF",
		X"2A",X"3A",X"80",X"50",X"0F",X"0F",X"0F",X"0F",X"E6",X"03",X"FE",X"03",X"20",X"08",X"06",X"2A",
		X"CD",X"DF",X"2A",X"C3",X"63",X"31",X"07",X"5F",X"D5",X"06",X"2B",X"CD",X"DF",X"2A",X"06",X"2E",
		X"CD",X"DF",X"2A",X"D1",X"16",X"00",X"21",X"7F",X"32",X"19",X"7E",X"32",X"2A",X"42",X"23",X"7E",
		X"32",X"4A",X"42",X"3A",X"80",X"50",X"0F",X"0F",X"E6",X"03",X"F6",X"02",X"C6",X"31",X"FE",X"34",
		X"20",X"01",X"3C",X"32",X"AC",X"41",X"06",X"29",X"CD",X"DF",X"2A",X"3A",X"40",X"50",X"07",X"E6",
		X"01",X"C6",X"2C",X"47",X"CD",X"DF",X"2A",X"3A",X"80",X"50",X"E6",X"08",X"CA",X"CF",X"30",X"AF",
		X"32",X"00",X"50",X"F3",X"21",X"07",X"50",X"AF",X"77",X"2D",X"20",X"FC",X"31",X"50",X"3A",X"06",
		X"03",X"D9",X"E1",X"D1",X"32",X"C0",X"50",X"C1",X"3E",X"3C",X"77",X"23",X"72",X"23",X"10",X"F8",
		X"3B",X"3B",X"C1",X"71",X"23",X"3E",X"3F",X"77",X"23",X"10",X"F8",X"3B",X"3B",X"1D",X"C2",X"A4",
		X"31",X"F1",X"D9",X"10",X"DC",X"31",X"C0",X"4F",X"06",X"30",X"CD",X"6D",X"32",X"10",X"FB",X"18",
		X"74",X"DD",X"E5",X"E5",X"AF",X"3E",X"40",X"C6",X"0C",X"67",X"3E",X"5A",X"C6",X"10",X"6F",X"E5",
		X"DD",X"E1",X"3E",X"50",X"DD",X"36",X"00",X"C0",X"DD",X"77",X"01",X"DD",X"36",X"02",X"80",X"DD",
		X"77",X"03",X"DD",X"36",X"04",X"C0",X"DD",X"77",X"05",X"E1",X"DD",X"E1",X"C9",X"32",X"C0",X"50",
		X"3A",X"40",X"50",X"E6",X"10",X"28",X"F6",X"3A",X"40",X"50",X"E6",X"27",X"C2",X"6C",X"00",X"06",
		X"08",X"CD",X"6D",X"32",X"10",X"FB",X"3A",X"40",X"50",X"E6",X"10",X"C2",X"6C",X"00",X"1E",X"01",
		X"06",X"04",X"32",X"C0",X"50",X"CD",X"6D",X"32",X"3A",X"00",X"50",X"A3",X"20",X"F4",X"CD",X"6D",
		X"32",X"32",X"C0",X"50",X"3A",X"00",X"50",X"EE",X"FF",X"20",X"F3",X"10",X"E5",X"CB",X"03",X"7B",
		X"FE",X"10",X"DA",X"20",X"32",X"21",X"00",X"40",X"06",X"04",X"3E",X"40",X"77",X"2C",X"20",X"FC",
		X"24",X"10",X"F7",X"00",X"00",X"00",X"3E",X"40",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F7",X"32",
		X"C0",X"50",X"3A",X"40",X"50",X"E6",X"10",X"CA",X"5F",X"32",X"C3",X"6C",X"00",X"32",X"C0",X"50",
		X"21",X"00",X"28",X"2B",X"7C",X"B5",X"20",X"FB",X"C9",X"CD",X"6D",X"32",X"10",X"FB",X"C9",X"30",
		X"32",X"30",X"34",X"30",X"38",X"00",X"FF",X"01",X"00",X"00",X"01",X"FF",X"00",X"00",X"FF",X"01",
		X"00",X"00",X"01",X"FF",X"00",X"00",X"FF",X"01",X"00",X"00",X"01",X"FF",X"00",X"00",X"FF",X"01",
		X"00",X"00",X"01",X"FF",X"00",X"55",X"2A",X"55",X"2A",X"55",X"55",X"55",X"55",X"55",X"2A",X"55",
		X"2A",X"52",X"4A",X"A5",X"94",X"25",X"25",X"25",X"25",X"22",X"22",X"22",X"22",X"01",X"01",X"01",
		X"01",X"58",X"02",X"08",X"07",X"60",X"09",X"10",X"0E",X"68",X"10",X"70",X"17",X"14",X"19",X"52",
		X"4A",X"A5",X"94",X"AA",X"2A",X"55",X"55",X"55",X"2A",X"55",X"2A",X"52",X"4A",X"A5",X"94",X"92",
		X"24",X"25",X"49",X"48",X"24",X"22",X"91",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"2A",X"55",X"2A",X"55",X"55",X"55",
		X"55",X"AA",X"2A",X"55",X"55",X"55",X"2A",X"55",X"2A",X"52",X"4A",X"A5",X"94",X"48",X"24",X"22",
		X"91",X"21",X"44",X"44",X"08",X"58",X"02",X"34",X"08",X"D8",X"09",X"B4",X"0F",X"58",X"11",X"08",
		X"16",X"34",X"17",X"55",X"55",X"55",X"55",X"D5",X"6A",X"D5",X"6A",X"AA",X"6A",X"55",X"D5",X"55",
		X"55",X"55",X"55",X"AA",X"2A",X"55",X"55",X"92",X"24",X"92",X"24",X"22",X"22",X"22",X"22",X"A4",
		X"01",X"54",X"06",X"F8",X"07",X"A8",X"0C",X"D4",X"0D",X"84",X"12",X"B0",X"13",X"D5",X"6A",X"D5",
		X"6A",X"D6",X"5A",X"AD",X"B5",X"D6",X"5A",X"AD",X"B5",X"D5",X"6A",X"D5",X"6A",X"AA",X"6A",X"55",
		X"D5",X"92",X"24",X"25",X"49",X"48",X"24",X"22",X"91",X"A4",X"01",X"54",X"06",X"F8",X"07",X"A8",
		X"0C",X"D4",X"0D",X"FE",X"FF",X"FF",X"FF",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"B6",
		X"6D",X"6D",X"DB",X"6D",X"6D",X"6D",X"6D",X"D6",X"5A",X"AD",X"B5",X"25",X"25",X"25",X"25",X"92",
		X"24",X"92",X"24",X"2C",X"01",X"DC",X"05",X"08",X"07",X"B8",X"0B",X"E4",X"0C",X"FE",X"FF",X"FF",
		X"FF",X"D5",X"6A",X"D5",X"6A",X"D5",X"6A",X"D5",X"6A",X"B6",X"6D",X"6D",X"DB",X"6D",X"6D",X"6D",
		X"6D",X"D6",X"5A",X"AD",X"B5",X"48",X"24",X"22",X"91",X"92",X"24",X"92",X"24",X"2C",X"01",X"DC",
		X"05",X"08",X"07",X"B8",X"0B",X"E4",X"0C",X"FE",X"FF",X"FF",X"FF",X"0E",X"00",X"C3",X"FD",X"33",
		X"0E",X"0C",X"C3",X"FD",X"33",X"0E",X"18",X"C3",X"FD",X"33",X"0E",X"24",X"C3",X"FD",X"33",X"0E",
		X"30",X"C3",X"FD",X"33",X"0E",X"3C",X"C3",X"FD",X"33",X"0E",X"48",X"C3",X"FD",X"33",X"0E",X"54",
		X"C3",X"FD",X"33",X"0E",X"60",X"C3",X"FD",X"33",X"0E",X"6C",X"C3",X"FD",X"33",X"3A",X"00",X"4F",
		X"A7",X"CC",X"7B",X"35",X"06",X"06",X"DD",X"21",X"0C",X"4F",X"DD",X"6E",X"00",X"DD",X"66",X"01",
		X"7E",X"FE",X"F0",X"CA",X"3F",X"34",X"FE",X"F1",X"CA",X"CC",X"34",X"FE",X"F2",X"CA",X"F8",X"34",
		X"FE",X"F3",X"CA",X"D8",X"34",X"FE",X"F5",X"CA",X"71",X"35",X"FE",X"F6",X"CA",X"05",X"35",X"FE",
		X"F7",X"CA",X"5D",X"35",X"FE",X"F8",X"CA",X"67",X"35",X"FE",X"FF",X"CA",X"2C",X"35",X"76",X"E5",
		X"3E",X"01",X"D7",X"4F",X"21",X"2E",X"4F",X"DF",X"79",X"84",X"CD",X"B7",X"34",X"12",X"CD",X"AB",
		X"35",X"DF",X"7C",X"81",X"12",X"E1",X"E5",X"3E",X"02",X"D7",X"4F",X"21",X"2E",X"4F",X"DF",X"79",
		X"85",X"CD",X"B7",X"34",X"1B",X"12",X"CD",X"AB",X"35",X"DF",X"7D",X"81",X"1B",X"12",X"21",X"0F",
		X"4F",X"78",X"D7",X"E5",X"3C",X"4F",X"21",X"3E",X"4F",X"DF",X"79",X"CB",X"2F",X"D7",X"FE",X"FF",
		X"C2",X"87",X"34",X"0E",X"00",X"18",X"EF",X"E1",X"71",X"5F",X"E1",X"3E",X"03",X"D7",X"57",X"D5",
		X"21",X"4E",X"4F",X"DF",X"E1",X"EB",X"72",X"2B",X"3A",X"09",X"4E",X"4F",X"3A",X"72",X"4E",X"A1",
		X"28",X"04",X"3E",X"C0",X"AB",X"5F",X"73",X"21",X"17",X"4F",X"78",X"D7",X"3D",X"77",X"11",X"00",
		X"00",X"20",X"62",X"1E",X"04",X"18",X"5E",X"4F",X"CB",X"29",X"CB",X"29",X"CB",X"29",X"CB",X"29",
		X"A7",X"F2",X"C9",X"34",X"F6",X"F0",X"0C",X"18",X"02",X"E6",X"0F",X"C9",X"EB",X"CD",X"AB",X"35",
		X"EB",X"D5",X"23",X"56",X"23",X"5E",X"18",X"13",X"EB",X"21",X"0F",X"4F",X"78",X"D7",X"36",X"00",
		X"EB",X"11",X"3E",X"4F",X"D5",X"23",X"5E",X"23",X"56",X"18",X"00",X"E1",X"D5",X"DF",X"EB",X"D1",
		X"72",X"2B",X"73",X"11",X"03",X"00",X"18",X"1D",X"23",X"4E",X"21",X"17",X"4F",X"78",X"D7",X"71",
		X"11",X"02",X"00",X"18",X"10",X"21",X"17",X"4F",X"78",X"D7",X"3D",X"77",X"11",X"00",X"00",X"20",
		X"04",X"1E",X"01",X"18",X"00",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"19",X"DD",X"75",X"00",X"DD",
		X"74",X"01",X"DD",X"2B",X"DD",X"2B",X"10",X"01",X"C9",X"C3",X"0A",X"34",X"21",X"1F",X"4F",X"78",
		X"D7",X"36",X"01",X"21",X"20",X"4F",X"7E",X"23",X"A6",X"23",X"A6",X"23",X"A6",X"23",X"A6",X"23",
		X"A6",X"11",X"00",X"00",X"28",X"CF",X"3A",X"02",X"4E",X"A7",X"CA",X"54",X"35",X"AF",X"32",X"00",
		X"4F",X"C3",X"8F",X"06",X"F7",X"45",X"00",X"00",X"21",X"04",X"4E",X"34",X"C9",X"78",X"EF",X"1C",
		X"30",X"47",X"11",X"01",X"00",X"18",X"AE",X"3E",X"40",X"32",X"AC",X"42",X"11",X"01",X"00",X"18",
		X"A4",X"23",X"7E",X"32",X"BC",X"4E",X"11",X"02",X"00",X"18",X"9A",X"3A",X"02",X"4E",X"A7",X"20",
		X"08",X"3E",X"02",X"32",X"CC",X"4E",X"32",X"DC",X"4E",X"21",X"2D",X"81",X"06",X"00",X"09",X"11",
		X"02",X"4F",X"01",X"0C",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"00",X"4F",X"32",X"A4",X"4D",X"21",
		X"1F",X"4F",X"3E",X"00",X"32",X"A5",X"4D",X"06",X"14",X"CF",X"C9",X"78",X"FE",X"06",X"20",X"04",
		X"21",X"C6",X"4D",X"C9",X"21",X"FE",X"4C",X"C9",X"05",X"C5",X"78",X"FE",X"01",X"28",X"04",X"06",
		X"00",X"18",X"06",X"3A",X"13",X"4E",X"E6",X"0F",X"47",X"DF",X"C1",X"C3",X"19",X"2C",X"CB",X"77",
		X"CA",X"30",X"1F",X"3E",X"01",X"02",X"C9",X"21",X"00",X"00",X"22",X"D2",X"4D",X"C9",X"3A",X"08",
		X"4D",X"E6",X"0F",X"CB",X"3F",X"CB",X"3F",X"2F",X"1E",X"1C",X"83",X"FE",X"18",X"20",X"02",X"3E",
		X"36",X"32",X"0A",X"4C",X"C9",X"03",X"04",X"01",X"02",X"01",X"01",X"01",X"01",X"0C",X"01",X"01",
		X"04",X"01",X"01",X"01",X"E8",X"4D",X"44",X"37",X"53",X"37",X"62",X"37",X"70",X"37",X"80",X"37",
		X"90",X"37",X"9C",X"37",X"B3",X"37",X"C7",X"37",X"B4",X"3C",X"93",X"3C",X"BE",X"B4",X"DA",X"B4",
		X"2C",X"3D",X"FF",X"3C",X"50",X"3D",X"16",X"38",X"24",X"38",X"CF",X"3C",X"D8",X"3C",X"22",X"3D",
		X"EF",X"3C",X"36",X"3D",X"01",X"00",X"02",X"00",X"03",X"00",X"66",X"38",X"6E",X"38",X"CE",X"3B",
		X"82",X"38",X"8C",X"38",X"96",X"38",X"A0",X"38",X"AA",X"38",X"B4",X"38",X"C4",X"38",X"19",X"39",
		X"D4",X"38",X"02",X"39",X"EB",X"38",X"6A",X"3D",X"30",X"39",X"41",X"39",X"5A",X"39",X"67",X"39",
		X"74",X"39",X"0D",X"3D",X"74",X"3D",X"1B",X"3D",X"8D",X"3D",X"06",X"3D",X"6A",X"3D",X"14",X"3D",
		X"83",X"3D",X"DE",X"37",X"D4",X"83",X"4D",X"49",X"4B",X"59",X"40",X"43",X"48",X"45",X"4C",X"4F",
		X"2F",X"81",X"2F",X"80",X"8C",X"02",X"4D",X"4D",X"4D",X"4D",X"4D",X"4D",X"4D",X"4D",X"4D",X"4D",
		X"2F",X"85",X"2F",X"80",X"8D",X"02",X"49",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"49",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"40",X"49",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"40",X"40",X"49",X"40",X"40",X"40",X"40",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"40",X"40",X"40",X"49",X"40",X"40",X"40",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"40",X"40",X"40",X"40",X"49",X"40",X"40",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"40",X"40",X"40",X"40",X"40",X"49",X"40",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"49",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"49",X"40",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"49",
		X"2F",X"89",X"2F",X"80",X"8D",X"02",X"49",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"2F",X"89",X"2F",X"80",X"3B",X"80",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"40",X"40",X"2F",
		X"8F",X"2F",X"80",X"3B",X"80",X"46",X"52",X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"2F",X"8F",
		X"2F",X"80",X"8C",X"02",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"45",X"2F",X"85",
		X"8C",X"02",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"54",X"57",X"4F",X"2F",X"85",X"2F",X"80",
		X"92",X"02",X"47",X"41",X"4D",X"45",X"40",X"40",X"4F",X"56",X"45",X"52",X"2F",X"81",X"2F",X"80",
		X"52",X"02",X"52",X"45",X"41",X"44",X"59",X"5B",X"2F",X"89",X"2F",X"90",X"ED",X"02",X"50",X"55",
		X"53",X"48",X"40",X"53",X"54",X"41",X"52",X"54",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"2F",
		X"87",X"2F",X"80",X"AF",X"02",X"31",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",
		X"4C",X"59",X"40",X"2F",X"87",X"2F",X"80",X"AF",X"02",X"31",X"40",X"4F",X"52",X"40",X"32",X"40",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"2F",X"87",X"00",X"2F",X"00",X"80",X"00",X"B1",X"02",
		X"32",X"40",X"4F",X"52",X"40",X"34",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"2F",X"87",
		X"00",X"2F",X"00",X"80",X"00",X"96",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"50",X"55",X"43",
		X"4B",X"4D",X"41",X"4E",X"40",X"46",X"4F",X"52",X"40",X"40",X"40",X"30",X"30",X"30",X"40",X"5D",
		X"5E",X"5F",X"2F",X"8E",X"2F",X"80",X"76",X"02",X"10",X"40",X"31",X"30",X"40",X"5D",X"5E",X"5F",
		X"2F",X"9F",X"2F",X"80",X"78",X"02",X"14",X"40",X"35",X"30",X"40",X"5D",X"5E",X"5F",X"2F",X"9F",
		X"2F",X"80",X"5D",X"02",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"83",X"2F",X"80",X"C5",
		X"02",X"40",X"2F",X"81",X"2F",X"80",X"C5",X"02",X"40",X"2F",X"81",X"2F",X"80",X"C8",X"02",X"40",
		X"2F",X"83",X"2F",X"80",X"C8",X"02",X"40",X"52",X"4F",X"4D",X"50",X"3B",X"3B",X"3B",X"3B",X"3B",
		X"3B",X"3B",X"2F",X"83",X"2F",X"80",X"25",X"80",X"81",X"85",X"2F",X"81",X"2F",X"90",X"6E",X"02",
		X"53",X"55",X"50",X"45",X"52",X"40",X"50",X"41",X"43",X"3B",X"4D",X"41",X"4E",X"2F",X"89",X"2F",
		X"80",X"4D",X"41",X"4E",X"2F",X"89",X"2F",X"80",X"2F",X"90",X"00",X"00",X"2E",X"80",X"86",X"8B",
		X"8D",X"8E",X"2F",X"8F",X"2F",X"90",X"30",X"80",X"40",X"40",X"40",X"40",X"2F",X"94",X"2F",X"90",
		X"32",X"80",X"89",X"8A",X"8D",X"8E",X"2F",X"89",X"2F",X"90",X"34",X"80",X"89",X"8A",X"8D",X"8E",
		X"2F",X"89",X"2F",X"90",X"04",X"03",X"4D",X"45",X"4D",X"4F",X"52",X"59",X"40",X"40",X"4F",X"4B",
		X"2F",X"8F",X"2F",X"80",X"04",X"03",X"42",X"41",X"44",X"40",X"40",X"40",X"40",X"52",X"40",X"4D",
		X"2F",X"8F",X"2F",X"80",X"08",X"03",X"31",X"40",X"43",X"4F",X"49",X"4E",X"40",X"40",X"31",X"40",
		X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"2F",X"8F",X"2F",X"80",X"08",X"03",X"32",X"40",X"43",
		X"4F",X"49",X"4E",X"53",X"40",X"31",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"2F",X"8F",
		X"2F",X"80",X"08",X"03",X"31",X"40",X"43",X"4F",X"49",X"4E",X"40",X"40",X"32",X"40",X"43",X"52",
		X"45",X"44",X"49",X"54",X"53",X"2F",X"8F",X"2F",X"80",X"08",X"03",X"46",X"52",X"45",X"45",X"40",
		X"40",X"50",X"4C",X"41",X"59",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"2F",X"8F",X"2F",X"80",
		X"0A",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"40",X"4E",X"4F",X"4E",X"45",X"2F",X"8F",X"2F",
		X"80",X"0A",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"2F",X"8F",X"2F",X"80",X"0C",X"03",X"50",
		X"55",X"43",X"4B",X"4D",X"41",X"4E",X"2F",X"8F",X"2F",X"80",X"0E",X"03",X"54",X"41",X"42",X"4C",
		X"45",X"40",X"40",X"2F",X"8F",X"2F",X"80",X"0E",X"03",X"55",X"50",X"52",X"49",X"47",X"48",X"54",
		X"2F",X"8F",X"2F",X"80",X"0A",X"02",X"30",X"30",X"30",X"2F",X"8F",X"2F",X"80",X"6B",X"01",X"40",
		X"2F",X"85",X"2F",X"3D",X"59",X"02",X"B6",X"02",X"C3",X"02",X"D0",X"02",X"C3",X"02",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"16",X"B5",X"25",X"B5",X"78",X"02",X"97",X"02",X"1F",X"03",
		X"3D",X"03",X"E6",X"02",X"06",X"B5",X"5B",X"03",X"6B",X"03",X"7B",X"03",X"8B",X"03",X"9B",X"03",
		X"AB",X"03",X"BB",X"03",X"CB",X"03",X"DB",X"03",X"EB",X"03",X"6A",X"B5",X"7A",X"B5",X"8A",X"B5",
		X"9A",X"B5",X"BA",X"B5",X"AA",X"B5",X"34",X"B5",X"43",X"B5",X"50",X"B5",X"5D",X"B5",X"AC",X"B4",
		X"94",X"36",X"A4",X"36",X"B4",X"36",X"C4",X"36",X"D4",X"36",X"E4",X"36",X"F4",X"36",X"04",X"37",
		X"14",X"37",X"24",X"37",X"34",X"37",X"04",X"1C",X"02",X"02",X"0A",X"01",X"11",X"02",X"02",X"0C",
		X"01",X"01",X"0E",X"01",X"01",X"01",X"01",X"03",X"01",X"07",X"1A",X"01",X"01",X"03",X"13",X"01",
		X"01",X"05",X"18",X"04",X"03",X"07",X"01",X"03",X"0E",X"04",X"0C",X"01",X"0F",X"01",X"01",X"01",
		X"01",X"04",X"02",X"07",X"16",X"02",X"02",X"03",X"01",X"01",X"01",X"01",X"0F",X"01",X"01",X"01",
		X"03",X"02",X"02",X"15",X"03",X"04",X"01",X"01",X"01",X"01",X"15",X"03",X"0B",X"01",X"01",X"01",
		X"01",X"0F",X"01",X"01",X"01",X"3C",X"01",X"01",X"01",X"01",X"0A",X"01",X"01",X"01",X"01",X"0F",
		X"0E",X"13",X"0E",X"11",X"0E",X"11",X"01",X"01",X"01",X"01",X"0A",X"01",X"01",X"01",X"01",X"00",
		X"02",X"40",X"01",X"3E",X"3D",X"10",X"40",X"40",X"0E",X"3D",X"3E",X"10",X"C2",X"43",X"01",X"3E",
		X"3D",X"10",X"21",X"C3",X"40",X"11",X"E6",X"39",X"36",X"14",X"1A",X"A7",X"C8",X"13",X"85",X"6F",
		X"D2",X"68",X"3A",X"24",X"18",X"F2",X"90",X"14",X"94",X"0F",X"98",X"15",X"9C",X"07",X"A0",X"14",
		X"A4",X"17",X"A8",X"16",X"AC",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"16",X"9C",X"16",X"9C",X"16",X"73",X"20",
		X"00",X"0C",X"00",X"0A",X"1F",X"00",X"72",X"20",X"FB",X"87",X"00",X"02",X"0F",X"00",X"59",X"01",
		X"06",X"08",X"00",X"00",X"02",X"00",X"59",X"01",X"06",X"09",X"00",X"00",X"02",X"00",X"59",X"02",
		X"06",X"0A",X"00",X"00",X"02",X"00",X"59",X"03",X"06",X"0B",X"00",X"00",X"02",X"00",X"59",X"04",
		X"06",X"0C",X"00",X"06",X"02",X"00",X"24",X"00",X"06",X"08",X"02",X"00",X"0A",X"00",X"36",X"07",
		X"87",X"6F",X"00",X"00",X"04",X"00",X"70",X"04",X"00",X"00",X"00",X"00",X"08",X"00",X"1C",X"70",
		X"8B",X"08",X"00",X"01",X"06",X"00",X"1C",X"70",X"8B",X"08",X"00",X"01",X"06",X"00",X"56",X"0C",
		X"FF",X"8C",X"00",X"02",X"08",X"00",X"56",X"00",X"02",X"0A",X"07",X"03",X"0C",X"00",X"36",X"38",
		X"FE",X"12",X"F8",X"04",X"0F",X"FC",X"22",X"01",X"01",X"06",X"00",X"01",X"07",X"00",X"01",X"02",
		X"04",X"08",X"10",X"20",X"40",X"80",X"01",X"03",X"06",X"0C",X"18",X"30",X"60",X"00",X"57",X"5C",
		X"61",X"67",X"6D",X"74",X"7B",X"82",X"8A",X"92",X"9A",X"A3",X"AD",X"B8",X"C3",X"D4",X"3B",X"F3",
		X"3B",X"58",X"3C",X"95",X"3C",X"DE",X"3C",X"DF",X"3C",X"01",X"02",X"01",X"1B",X"03",X"03",X"1A",
		X"03",X"03",X"1A",X"03",X"03",X"1A",X"01",X"01",X"01",X"01",X"01",X"01",X"5A",X"01",X"01",X"01",
		X"01",X"01",X"21",X"20",X"20",X"1A",X"01",X"01",X"01",X"01",X"01",X"61",X"20",X"20",X"20",X"1A",
		X"01",X"01",X"01",X"01",X"01",X"01",X"5B",X"04",X"1B",X"06",X"1A",X"06",X"1A",X"06",X"1B",X"01",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"06",X"1A",X"06",X"1A",X"06",X"1B",X"01",X"01",
		X"01",X"F1",X"03",X"F2",X"03",X"F3",X"0A",X"F4",X"02",X"90",X"7C",X"7B",X"7A",X"79",X"79",X"78",
		X"97",X"76",X"75",X"74",X"73",X"72",X"91",X"A8",X"88",X"60",X"4A",X"4C",X"91",X"95",X"88",X"95",
		X"91",X"95",X"88",X"95",X"91",X"95",X"88",X"95",X"95",X"98",X"94",X"97",X"93",X"96",X"88",X"96",
		X"93",X"96",X"88",X"96",X"93",X"96",X"88",X"96",X"B6",X"B3",X"75",X"76",X"77",X"78",X"78",X"75",
		X"73",X"68",X"91",X"95",X"88",X"95",X"91",X"95",X"88",X"95",X"86",X"96",X"95",X"92",X"93",X"8C",
		X"8A",X"88",X"86",X"90",X"90",X"96",X"95",X"90",X"90",X"86",X"90",X"96",X"90",X"96",X"91",X"88",
		X"81",X"FF",X"47",X"30",X"4B",X"10",X"4C",X"10",X"4D",X"10",X"4E",X"10",X"77",X"20",X"4E",X"10",
		X"4D",X"10",X"4C",X"10",X"4A",X"10",X"47",X"10",X"46",X"10",X"65",X"30",X"66",X"30",X"67",X"40",
		X"70",X"F0",X"FB",X"3B",X"F1",X"00",X"F2",X"02",X"F3",X"0A",X"F4",X"00",X"88",X"6C",X"71",X"72",
		X"73",X"73",X"71",X"93",X"6C",X"73",X"75",X"76",X"76",X"75",X"96",X"7C",X"7A",X"78",X"76",X"75",
		X"96",X"6C",X"91",X"A0",X"88",X"75",X"76",X"77",X"78",X"71",X"73",X"74",X"75",X"71",X"75",X"71",
		X"68",X"68",X"65",X"66",X"67",X"A8",X"AB",X"AC",X"8C",X"86",X"76",X"75",X"6C",X"71",X"75",X"73",
		X"6B",X"6C",X"73",X"76",X"7A",X"78",X"78",X"76",X"73",X"6C",X"AA",X"A8",X"71",X"73",X"74",X"75",
		X"6A",X"6B",X"6C",X"73",X"75",X"76",X"77",X"78",X"71",X"73",X"74",X"75",X"71",X"75",X"71",X"68",
		X"48",X"40",X"68",X"67",X"68",X"AA",X"A9",X"AA",X"6A",X"60",X"8A",X"76",X"75",X"73",X"71",X"71",
		X"73",X"95",X"75",X"73",X"71",X"68",X"68",X"61",X"63",X"6A",X"A8",X"6C",X"76",X"6A",X"6C",X"91",
		X"90",X"91",X"FF",X"96",X"03",X"40",X"41",X"44",X"44",X"49",X"54",X"49",X"4F",X"4E",X"41",X"4C",
		X"40",X"40",X"40",X"40",X"41",X"54",X"40",X"40",X"40",X"30",X"30",X"30",X"40",X"5D",X"5E",X"5F",
		X"2F",X"95",X"2F",X"80",X"5A",X"02",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"2F",X"07",X"07",
		X"07",X"01",X"01",X"01",X"01",X"2F",X"80",X"50",X"40",X"40",X"40",X"2F",X"87",X"2F",X"80",X"5B",
		X"02",X"40",X"2F",X"81",X"2F",X"80",X"2F",X"80",X"92",X"02",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"2F",X"81",X"2F",X"80",X"6E",X"02",X"40",X"2F",X"81",X"2F",X"80",X"92",
		X"02",X"40",X"40",X"54",X"55",X"52",X"42",X"4F",X"5B",X"40",X"40",X"2F",X"89",X"2F",X"80",X"6E",
		X"02",X"40",X"2F",X"83",X"2F",X"80",X"6E",X"02",X"40",X"2F",X"89",X"2F",X"80",X"6E",X"02",X"40",
		X"2F",X"85",X"2F",X"80",X"3D",X"02",X"40",X"2F",X"81",X"2F",X"80",X"6E",X"02",X"40",X"2F",X"87",
		X"2F",X"80",X"2F",X"02",X"4D",X"49",X"4B",X"59",X"2F",X"87",X"2F",X"80",X"2F",X"02",X"4D",X"49",
		X"4B",X"59",X"2F",X"85",X"2F",X"80",X"49",X"03",X"41",X"54",X"52",X"41",X"50",X"41",X"4E",X"44",
		X"4F",X"40",X"55",X"4E",X"40",X"43",X"4F",X"52",X"41",X"5A",X"4F",X"4E",X"2F",X"88",X"2F",X"80",
		X"53",X"03",X"56",X"49",X"44",X"41",X"40",X"45",X"58",X"54",X"52",X"41",X"40",X"4F",X"40",X"50",
		X"55",X"4E",X"54",X"41",X"47",X"45",X"2F",X"82",X"2F",X"80",X"2F",X"02",X"40",X"40",X"40",X"40",
		X"2F",X"8F",X"2F",X"80",X"6B",X"02",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"2F",
		X"85",X"2F",X"80",X"2F",X"02",X"40",X"40",X"40",X"40",X"2F",X"87",X"2F",X"80",X"6B",X"02",X"40",
		X"2F",X"8F",X"2F",X"80",X"0C",X"03",X"40",X"2F",X"8F",X"2F",X"80",X"3A",X"78",X"4C",X"E6",X"0F",
		X"E7",X"6A",X"3E",X"C1",X"3D",X"D9",X"3E",X"76",X"80",X"BC",X"80",X"FA",X"80",X"BC",X"80",X"91",
		X"80",X"C9",X"3D",X"D9",X"3E",X"9F",X"80",X"FA",X"80",X"C9",X"3D",X"BC",X"80",X"83",X"80",X"FA",
		X"80",X"3E",X"02",X"32",X"70",X"4C",X"C3",X"C9",X"3D",X"3A",X"02",X"4E",X"FE",X"10",X"C4",X"04",
		X"97",X"3A",X"02",X"4E",X"E7",X"CA",X"B5",X"F8",X"3D",X"FE",X"3D",X"0C",X"00",X"CB",X"33",X"04",
		X"3E",X"D0",X"33",X"0A",X"3E",X"D5",X"33",X"10",X"3E",X"DA",X"33",X"1C",X"3E",X"DF",X"33",X"1C",
		X"3E",X"1C",X"3E",X"1C",X"3E",X"08",X"3F",X"C9",X"EF",X"20",X"21",X"C3",X"8F",X"06",X"EF",X"20",
		X"1B",X"C3",X"8F",X"06",X"EF",X"20",X"1C",X"C3",X"8F",X"06",X"EF",X"20",X"1D",X"C3",X"8F",X"06",
		X"EF",X"20",X"1E",X"C3",X"8F",X"06",X"EF",X"20",X"1F",X"C3",X"8F",X"06",X"EF",X"20",X"20",X"C3",
		X"8F",X"06",X"EF",X"20",X"22",X"C3",X"8F",X"06",X"EF",X"20",X"23",X"C3",X"8F",X"06",X"EF",X"20",
		X"24",X"C3",X"8F",X"06",X"3A",X"01",X"4F",X"E6",X"10",X"20",X"0A",X"EF",X"1C",X"0C",X"EF",X"20",
		X"0A",X"EF",X"20",X"25",X"C9",X"EF",X"1C",X"0D",X"EF",X"20",X"09",X"C9",X"3A",X"01",X"4F",X"E6",
		X"10",X"20",X"07",X"EF",X"20",X"0A",X"EF",X"20",X"25",X"C9",X"3E",X"99",X"CD",X"2C",X"AF",X"E6",
		X"01",X"28",X"F7",X"EF",X"20",X"09",X"C9",X"C3",X"8F",X"06",X"3A",X"02",X"4E",X"FE",X"00",X"20",
		X"68",X"3A",X"78",X"4C",X"A7",X"20",X"62",X"EF",X"30",X"25",X"3A",X"02",X"4E",X"FE",X"20",X"28",
		X"05",X"FE",X"10",X"D4",X"1B",X"97",X"E7",X"CA",X"B5",X"32",X"97",X"32",X"97",X"32",X"97",X"32",
		X"97",X"32",X"97",X"32",X"97",X"32",X"97",X"32",X"97",X"32",X"97",X"32",X"97",X"32",X"97",X"32",
		X"97",X"32",X"97",X"32",X"97",X"32",X"97",X"CA",X"B5",X"F8",X"3D",X"FE",X"3D",X"0C",X"00",X"CB",
		X"33",X"04",X"3E",X"D0",X"33",X"0A",X"3E",X"D5",X"33",X"10",X"3E",X"DA",X"33",X"1C",X"3E",X"DF",
		X"33",X"1C",X"3E",X"1C",X"3E",X"1C",X"3E",X"08",X"3F",X"C9",X"3A",X"01",X"4F",X"3C",X"E6",X"1F",
		X"32",X"01",X"4F",X"E6",X"0F",X"C0",X"C3",X"8F",X"06",X"3A",X"02",X"4E",X"FE",X"10",X"C4",X"1B",
		X"97",X"3A",X"02",X"4E",X"E7",X"CA",X"B5",X"F8",X"3D",X"FE",X"3D",X"0C",X"00",X"CB",X"33",X"04",
		X"3E",X"D0",X"33",X"0A",X"3E",X"D5",X"33",X"10",X"3E",X"DA",X"33",X"1C",X"3E",X"DF",X"33",X"1C",
		X"3E",X"1C",X"3E",X"1C",X"3E",X"08",X"3F",X"C9",X"AF",X"32",X"14",X"4E",X"3A",X"78",X"4C",X"E6",
		X"0F",X"32",X"13",X"4E",X"C3",X"82",X"06",X"3A",X"01",X"4F",X"3C",X"E6",X"1F",X"32",X"01",X"4F",
		X"E6",X"07",X"CD",X"2C",X"AF",X"E6",X"0F",X"E7",X"92",X"3F",X"38",X"3F",X"56",X"3F",X"74",X"3F",
		X"74",X"3F",X"56",X"3F",X"38",X"3F",X"92",X"3F",X"21",X"63",X"40",X"11",X"49",X"3B",X"36",X"10",
		X"7C",X"C6",X"04",X"67",X"36",X"01",X"7C",X"C6",X"FC",X"67",X"1A",X"A7",X"C8",X"13",X"85",X"6F",
		X"D2",X"3E",X"3F",X"24",X"18",X"E8",X"21",X"63",X"40",X"11",X"49",X"3B",X"36",X"12",X"7C",X"C6",
		X"04",X"67",X"36",X"07",X"7C",X"C6",X"FC",X"67",X"1A",X"A7",X"C8",X"13",X"85",X"6F",X"D2",X"5C",
		X"3F",X"24",X"18",X"E8",X"21",X"63",X"40",X"11",X"49",X"3B",X"36",X"14",X"7C",X"C6",X"04",X"67",
		X"36",X"0F",X"7C",X"C6",X"FC",X"67",X"1A",X"A7",X"C8",X"13",X"85",X"6F",X"D2",X"7A",X"3F",X"24",
		X"18",X"E8",X"21",X"63",X"40",X"11",X"49",X"3B",X"36",X"40",X"1A",X"A7",X"C8",X"13",X"85",X"6F",
		X"D2",X"98",X"3F",X"24",X"18",X"F2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AB",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"C5",X"E5",X"CD",X"A0",X"B3",X"E1",X"C1",X"F1");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
