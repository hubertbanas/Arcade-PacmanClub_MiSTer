library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C9",X"E6",X"07",X"CD",X"2C",X"AF",X"E6",X"00",X"E7",X"17",X"80",X"56",X"3F",X"74",X"3F",X"74",
		X"3F",X"56",X"3F",X"38",X"3F",X"92",X"3F",X"26",X"40",X"3A",X"01",X"4F",X"E6",X"0F",X"F6",X"60",
		X"C6",X"03",X"6F",X"2D",X"11",X"49",X"3B",X"36",X"40",X"7C",X"C6",X"04",X"67",X"36",X"0F",X"7C",
		X"C6",X"FC",X"67",X"1A",X"A7",X"28",X"09",X"13",X"85",X"6F",X"D2",X"27",X"80",X"24",X"18",X"E7",
		X"26",X"40",X"3A",X"01",X"4F",X"E6",X"0F",X"F6",X"60",X"C6",X"03",X"6F",X"11",X"49",X"3B",X"36",
		X"14",X"7C",X"C6",X"04",X"67",X"36",X"0F",X"7C",X"C6",X"FC",X"67",X"1A",X"A7",X"C8",X"13",X"85",
		X"6F",X"D2",X"4F",X"80",X"24",X"18",X"E8",X"C9",X"3E",X"00",X"32",X"70",X"4C",X"3E",X"01",X"32",
		X"13",X"4E",X"C3",X"08",X"3F",X"C9",X"3E",X"01",X"32",X"70",X"4C",X"3E",X"02",X"32",X"13",X"4E",
		X"C3",X"08",X"3F",X"3E",X"02",X"32",X"70",X"4C",X"3E",X"03",X"32",X"13",X"4E",X"C3",X"08",X"3F",
		X"C9",X"3E",X"01",X"32",X"70",X"4C",X"3E",X"09",X"32",X"13",X"4E",X"C3",X"08",X"3F",X"C9",X"3E",
		X"02",X"32",X"70",X"4C",X"3E",X"0C",X"32",X"13",X"4E",X"C3",X"08",X"3F",X"C9",X"3E",X"02",X"32",
		X"70",X"4C",X"3E",X"0D",X"32",X"13",X"4E",X"C3",X"08",X"3F",X"C9",X"C9",X"3A",X"02",X"4E",X"FE",
		X"18",X"C4",X"04",X"97",X"3A",X"02",X"4E",X"E7",X"CA",X"B5",X"F8",X"3D",X"FE",X"3D",X"0C",X"00",
		X"04",X"3E",X"0A",X"3E",X"10",X"3E",X"EE",X"33",X"10",X"3E",X"22",X"3E",X"F3",X"33",X"F8",X"33",
		X"2E",X"3E",X"FE",X"3D",X"FE",X"3D",X"04",X"3E",X"0A",X"3E",X"10",X"3E",X"10",X"3E",X"E4",X"33",
		X"22",X"3E",X"E9",X"33",X"1C",X"3E",X"DF",X"33",X"08",X"3F",X"AF",X"32",X"70",X"4C",X"3A",X"02",
		X"4E",X"FE",X"10",X"C4",X"04",X"97",X"3A",X"02",X"4E",X"E7",X"CA",X"B5",X"F8",X"3D",X"FE",X"3D",
		X"0C",X"00",X"CB",X"33",X"04",X"3E",X"D0",X"33",X"0A",X"3E",X"D5",X"33",X"10",X"3E",X"DA",X"33",
		X"E4",X"33",X"22",X"3E",X"E9",X"33",X"1C",X"3E",X"DF",X"33",X"08",X"3F",X"C9",X"42",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"65",X"82",X"75",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"65",X"82",X"98",X"82",X"A8",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"65",X"82",X"98",X"82",X"CB",X"82",X"EB",X"82",X"41",X"82",X"41",X"82",X"65",X"82",X"98",
		X"82",X"CB",X"82",X"FE",X"82",X"0E",X"83",X"41",X"82",X"65",X"82",X"98",X"82",X"CB",X"82",X"FE",
		X"82",X"41",X"82",X"2D",X"83",X"57",X"84",X"61",X"84",X"6B",X"84",X"75",X"84",X"41",X"82",X"43",
		X"83",X"42",X"82",X"75",X"82",X"A8",X"82",X"EB",X"82",X"41",X"82",X"89",X"83",X"57",X"84",X"61",
		X"84",X"6B",X"84",X"75",X"84",X"41",X"82",X"7F",X"84",X"55",X"82",X"88",X"82",X"BB",X"82",X"DB",
		X"82",X"0E",X"83",X"A5",X"83",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",X"82",X"41",
		X"82",X"FF",X"F1",X"00",X"80",X"F3",X"0A",X"84",X"F2",X"70",X"F0",X"10",X"00",X"01",X"F2",X"40",
		X"F0",X"10",X"00",X"01",X"FF",X"F3",X"0A",X"84",X"F2",X"70",X"F0",X"F0",X"00",X"01",X"F2",X"70",
		X"F0",X"10",X"00",X"01",X"FF",X"F3",X"0A",X"84",X"F2",X"70",X"F0",X"00",X"00",X"01",X"F2",X"40",
		X"F0",X"00",X"00",X"01",X"FF",X"F1",X"00",X"90",X"F3",X"0A",X"84",X"F2",X"70",X"F0",X"10",X"00",
		X"03",X"F2",X"40",X"F0",X"10",X"00",X"03",X"FF",X"F3",X"0A",X"84",X"F2",X"70",X"F0",X"F0",X"00",
		X"03",X"F2",X"70",X"F0",X"10",X"00",X"03",X"FF",X"F3",X"0A",X"84",X"F2",X"70",X"F0",X"00",X"00",
		X"03",X"F2",X"40",X"F0",X"00",X"00",X"03",X"FF",X"F1",X"00",X"A0",X"F3",X"0A",X"84",X"F2",X"70",
		X"F0",X"10",X"00",X"05",X"F2",X"40",X"F0",X"10",X"00",X"05",X"FF",X"F3",X"0A",X"84",X"F2",X"70",
		X"F0",X"F0",X"00",X"05",X"F2",X"70",X"F0",X"10",X"00",X"05",X"FF",X"F3",X"0A",X"84",X"F2",X"70",
		X"F0",X"00",X"00",X"05",X"F2",X"40",X"F0",X"00",X"00",X"05",X"FF",X"F3",X"0A",X"84",X"F2",X"70",
		X"F0",X"F0",X"00",X"07",X"F2",X"70",X"F0",X"10",X"00",X"07",X"FF",X"F1",X"00",X"B0",X"F3",X"0A",
		X"84",X"F2",X"70",X"F0",X"10",X"00",X"07",X"F2",X"40",X"F0",X"10",X"00",X"07",X"FF",X"F3",X"0A",
		X"84",X"F2",X"70",X"F0",X"00",X"00",X"07",X"F2",X"40",X"F0",X"00",X"00",X"07",X"FF",X"F1",X"00",
		X"C0",X"F3",X"E2",X"83",X"F2",X"70",X"F0",X"10",X"00",X"09",X"F2",X"40",X"F0",X"10",X"00",X"09",
		X"F2",X"70",X"F0",X"00",X"00",X"09",X"F2",X"40",X"F0",X"00",X"00",X"09",X"FF",X"F1",X"00",X"70",
		X"F3",X"D9",X"83",X"F2",X"40",X"F0",X"F0",X"00",X"05",X"F2",X"04",X"F3",X"EB",X"83",X"F0",X"00",
		X"10",X"05",X"FF",X"F2",X"01",X"F3",X"D9",X"83",X"F0",X"00",X"01",X"05",X"FF",X"06",X"40",X"0E",
		X"00",X"DD",X"21",X"00",X"00",X"DD",X"E5",X"E1",X"16",X"00",X"7E",X"5F",X"DD",X"19",X"E5",X"2A",
		X"6A",X"4C",X"77",X"E1",X"23",X"0B",X"79",X"B0",X"20",X"EE",X"11",X"00",X"40",X"19",X"01",X"00",
		X"40",X"16",X"00",X"7E",X"5F",X"DD",X"19",X"E5",X"2A",X"6A",X"4C",X"77",X"E1",X"23",X"0B",X"79",
		X"B0",X"20",X"EE",X"DD",X"E5",X"E1",X"7D",X"AF",X"C9",X"F1",X"00",X"90",X"F2",X"30",X"F3",X"E2",
		X"83",X"F0",X"00",X"00",X"05",X"F3",X"E2",X"83",X"F2",X"70",X"F0",X"10",X"00",X"05",X"F2",X"30",
		X"F0",X"10",X"00",X"05",X"FF",X"F3",X"D9",X"83",X"F2",X"70",X"F0",X"F0",X"00",X"05",X"F2",X"30",
		X"F0",X"F0",X"00",X"05",X"FF",X"1B",X"1B",X"19",X"19",X"1B",X"1B",X"32",X"32",X"FF",X"9B",X"9B",
		X"99",X"99",X"9B",X"9B",X"B2",X"B2",X"FF",X"6E",X"6E",X"5A",X"5A",X"6E",X"6E",X"72",X"72",X"FF",
		X"EE",X"EE",X"DA",X"DA",X"EE",X"EE",X"F2",X"F2",X"FF",X"37",X"37",X"2D",X"2D",X"37",X"37",X"2F",
		X"2F",X"FF",X"B7",X"B7",X"AD",X"AD",X"B7",X"B7",X"AF",X"AF",X"FF",X"36",X"36",X"F1",X"F1",X"36",
		X"36",X"F3",X"F3",X"FF",X"34",X"34",X"31",X"31",X"34",X"34",X"33",X"33",X"FF",X"24",X"24",X"24",
		X"25",X"25",X"25",X"A4",X"A4",X"A4",X"A5",X"A5",X"A5",X"FF",X"24",X"24",X"24",X"25",X"25",X"25",
		X"A4",X"A4",X"A4",X"A5",X"A5",X"A5",X"FF",X"26",X"26",X"26",X"27",X"27",X"27",X"FF",X"1F",X"FF",
		X"1E",X"FF",X"10",X"10",X"10",X"14",X"14",X"14",X"16",X"16",X"16",X"FF",X"11",X"11",X"11",X"15",
		X"15",X"15",X"17",X"17",X"17",X"FF",X"12",X"FF",X"13",X"FF",X"30",X"FF",X"18",X"18",X"18",X"18",
		X"2C",X"2C",X"2C",X"2C",X"FF",X"07",X"FF",X"0F",X"FF",X"00",X"FF",X"01",X"FF",X"02",X"FF",X"03",
		X"FF",X"04",X"FF",X"05",X"FF",X"06",X"FF",X"F3",X"FD",X"83",X"F0",X"E0",X"20",X"01",X"F2",X"50",
		X"FF",X"F3",X"FD",X"83",X"F0",X"20",X"20",X"03",X"F2",X"50",X"FF",X"F3",X"FD",X"83",X"F0",X"E0",
		X"E0",X"05",X"F2",X"50",X"FF",X"F3",X"FD",X"83",X"F0",X"20",X"E0",X"05",X"F2",X"50",X"FF",X"F3",
		X"E2",X"83",X"F0",X"00",X"00",X"09",X"F2",X"50",X"FF",X"F2",X"01",X"F3",X"55",X"84",X"F0",X"00",
		X"00",X"16",X"F2",X"01",X"F6",X"F2",X"01",X"FF",X"F2",X"01",X"F3",X"55",X"84",X"F0",X"00",X"00",
		X"16",X"F2",X"01",X"F6",X"F2",X"01",X"FF",X"F2",X"01",X"F3",X"4F",X"84",X"F0",X"00",X"00",X"07",
		X"F2",X"01",X"F6",X"F2",X"01",X"FF",X"F2",X"01",X"F3",X"55",X"84",X"F0",X"00",X"00",X"16",X"F2",
		X"01",X"F6",X"F2",X"01",X"FF",X"F2",X"01",X"F3",X"55",X"84",X"F0",X"00",X"00",X"16",X"F2",X"01",
		X"F6",X"F2",X"01",X"FF",X"F2",X"01",X"F3",X"55",X"84",X"F0",X"00",X"00",X"16",X"F2",X"01",X"F6",
		X"F2",X"01",X"FF",X"F2",X"01",X"F3",X"55",X"84",X"F0",X"00",X"00",X"16",X"F2",X"01",X"F6",X"F2",
		X"01",X"FF",X"F1",X"00",X"94",X"F3",X"B5",X"83",X"F2",X"72",X"F0",X"F0",X"00",X"09",X"F2",X"5F",
		X"F6",X"FF",X"F1",X"00",X"94",X"F3",X"B5",X"83",X"F2",X"72",X"F0",X"F0",X"00",X"09",X"F2",X"5F",
		X"F3",X"BE",X"83",X"F2",X"72",X"F0",X"14",X"00",X"09",X"F2",X"20",X"F6",X"FF",X"3A",X"09",X"4D",
		X"E6",X"07",X"CB",X"3F",X"2F",X"1E",X"30",X"83",X"CB",X"47",X"20",X"02",X"3E",X"37",X"32",X"0A",
		X"4C",X"C9",X"3A",X"08",X"4D",X"E6",X"07",X"CB",X"3F",X"1E",X"30",X"83",X"CB",X"47",X"20",X"02",
		X"3E",X"34",X"32",X"0A",X"4C",X"C9",X"3A",X"09",X"4D",X"E6",X"07",X"CB",X"3F",X"1E",X"AC",X"83",
		X"CB",X"47",X"20",X"02",X"3E",X"35",X"32",X"0A",X"4C",X"C9",X"3A",X"08",X"4D",X"E6",X"07",X"CB",
		X"3F",X"2F",X"1E",X"F4",X"83",X"CB",X"47",X"20",X"02",X"3E",X"36",X"32",X"0A",X"4C",X"C9",X"3A",
		X"0C",X"4C",X"FE",X"1E",X"C0",X"2A",X"26",X"4D",X"C9",X"3A",X"A4",X"4D",X"A7",X"C0",X"3A",X"D4",
		X"4D",X"A7",X"CA",X"D2",X"85",X"3A",X"D2",X"4D",X"A7",X"CA",X"D2",X"85",X"3A",X"41",X"4C",X"47",
		X"21",X"4C",X"87",X"DF",X"ED",X"5B",X"D2",X"4D",X"19",X"22",X"D2",X"4D",X"21",X"41",X"4C",X"34",
		X"7E",X"E6",X"0F",X"C0",X"21",X"40",X"4C",X"35",X"FA",X"68",X"86",X"7E",X"57",X"CB",X"3F",X"CB",
		X"3F",X"21",X"BC",X"4E",X"CB",X"EE",X"2A",X"42",X"4C",X"D7",X"4F",X"3E",X"03",X"A2",X"28",X"07",
		X"CB",X"39",X"CB",X"39",X"3D",X"20",X"F9",X"3E",X"03",X"A1",X"07",X"07",X"07",X"07",X"32",X"41",
		X"4C",X"C9",X"3A",X"70",X"4C",X"FE",X"02",X"20",X"1B",X"3A",X"0E",X"4E",X"FE",X"20",X"CA",X"05",
		X"86",X"FE",X"40",X"CA",X"05",X"86",X"FE",X"A0",X"CA",X"05",X"86",X"FE",X"D0",X"C0",X"21",X"0D",
		X"4E",X"C3",X"08",X"86",X"3A",X"0E",X"4E",X"FE",X"40",X"CA",X"05",X"86",X"FE",X"B0",X"C0",X"21",
		X"0D",X"4E",X"C3",X"08",X"86",X"21",X"0C",X"4E",X"7E",X"A7",X"C0",X"34",X"3A",X"13",X"4E",X"FE",
		X"07",X"38",X"0A",X"06",X"07",X"ED",X"5F",X"E6",X"1F",X"90",X"30",X"FD",X"80",X"21",X"50",X"86",
		X"47",X"87",X"80",X"D7",X"32",X"0C",X"4C",X"23",X"7E",X"32",X"0D",X"4C",X"23",X"7E",X"32",X"D4",
		X"4D",X"21",X"AB",X"86",X"CD",X"80",X"86",X"23",X"5E",X"23",X"56",X"ED",X"53",X"D2",X"4D",X"C9",
		X"00",X"14",X"01",X"0F",X"02",X"15",X"03",X"07",X"04",X"14",X"05",X"17",X"06",X"16",X"00",X"14",
		X"00",X"14",X"06",X"01",X"0F",X"07",X"02",X"15",X"08",X"00",X"14",X"09",X"04",X"14",X"0A",X"05",
		X"15",X"0B",X"06",X"16",X"0C",X"07",X"09",X"0D",X"3A",X"D3",X"4D",X"C6",X"20",X"FE",X"40",X"38",
		X"52",X"2A",X"42",X"4C",X"11",X"BB",X"86",X"37",X"3F",X"ED",X"52",X"20",X"23",X"21",X"B3",X"86",
		X"CD",X"A1",X"94",X"69",X"60",X"ED",X"5F",X"E6",X"03",X"47",X"87",X"87",X"80",X"D7",X"5F",X"23",
		X"56",X"ED",X"53",X"42",X"4C",X"23",X"7E",X"32",X"40",X"4C",X"3E",X"1F",X"32",X"41",X"4C",X"C9",
		X"21",X"BB",X"86",X"22",X"42",X"4C",X"3E",X"1D",X"C3",X"97",X"86",X"62",X"8A",X"5B",X"8D",X"3D",
		X"90",X"AC",X"93",X"95",X"8A",X"8E",X"8D",X"65",X"90",X"DF",X"93",X"FA",X"FF",X"55",X"55",X"01",
		X"80",X"AA",X"02",X"3A",X"70",X"4C",X"FE",X"03",X"CA",X"AF",X"11",X"3E",X"00",X"32",X"0D",X"4C",
		X"C3",X"AF",X"11",X"F5",X"ED",X"5B",X"D2",X"4D",X"7C",X"92",X"C6",X"03",X"FE",X"06",X"30",X"68",
		X"7D",X"93",X"C6",X"03",X"FE",X"06",X"30",X"60",X"3A",X"0C",X"4C",X"FE",X"1E",X"CD",X"15",X"87",
		X"3E",X"01",X"32",X"0D",X"4C",X"F1",X"C6",X"02",X"32",X"0C",X"4C",X"D6",X"02",X"C3",X"40",X"1C",
		X"3A",X"70",X"4C",X"FE",X"02",X"28",X"03",X"FE",X"03",X"C0",X"3A",X"14",X"4E",X"FE",X"06",X"D0",
		X"CD",X"BB",X"29",X"AF",X"C9",X"F5",X"DD",X"E5",X"3A",X"70",X"4C",X"FE",X"03",X"28",X"04",X"FE",
		X"02",X"20",X"21",X"3A",X"70",X"4C",X"FE",X"03",X"20",X"03",X"3E",X"40",X"77",X"CD",X"65",X"1D",
		X"DD",X"21",X"0D",X"42",X"DD",X"36",X"00",X"40",X"DD",X"36",X"01",X"40",X"DD",X"36",X"E0",X"40",
		X"DD",X"36",X"E1",X"40",X"DD",X"E1",X"F1",X"C9",X"F1",X"C3",X"52",X"1C",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"FF",X"FE",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"FE",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"01",X"FF",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"40",X"FC",X"D0",X"D2",
		X"D2",X"D2",X"D2",X"D4",X"FC",X"DA",X"02",X"DC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"DA",X"02",
		X"DC",X"DC",X"FC",X"FC",X"D0",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D4",X"FC",X"DA",X"05",
		X"DC",X"FC",X"DA",X"02",X"DC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"DA",X"02",X"DC",X"FC",X"FC",
		X"FC",X"DA",X"08",X"DC",X"FC",X"DA",X"02",X"E6",X"EA",X"02",X"E7",X"D2",X"EB",X"02",X"E7",X"D2",
		X"D2",X"D2",X"D2",X"D2",X"D2",X"EB",X"02",X"E7",X"D2",X"D2",X"D2",X"EB",X"02",X"E6",X"E8",X"E8",
		X"E8",X"EA",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"15",X"DE",X"C0",X"C0",X"C0",X"E4",X"02",
		X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"E6",X"E8",
		X"E8",X"E8",X"EA",X"02",X"E6",X"EA",X"02",X"E6",X"EA",X"02",X"DE",X"C0",X"C0",X"C0",X"E4",X"02",
		X"DC",X"FC",X"DA",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"F5",X"E4",X"02",X"DE",X"F3",
		X"E9",X"E9",X"EB",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"E7",X"E9",X"E9",X"E9",X"EB",X"02",
		X"DC",X"FC",X"DA",X"09",X"DE",X"E4",X"02",X"DE",X"E4",X"05",X"DE",X"E4",X"02",X"DE",X"E4",X"08",
		X"DC",X"FC",X"FA",X"E8",X"E8",X"EA",X"02",X"E6",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",
		X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"E8",X"EA",X"02",
		X"DC",X"FC",X"FB",X"E9",X"E9",X"EB",X"02",X"DE",X"C0",X"E4",X"02",X"E7",X"EB",X"02",X"E7",X"EB",
		X"02",X"E7",X"E9",X"E9",X"F5",X"E4",X"02",X"E7",X"EB",X"02",X"DE",X"F3",X"E9",X"E9",X"EB",X"02",
		X"DC",X"FC",X"DA",X"05",X"DE",X"C0",X"E4",X"0B",X"DE",X"E4",X"05",X"DE",X"E4",X"05",X"DC",X"FC",
		X"DA",X"02",X"E6",X"EA",X"02",X"DE",X"C0",X"E4",X"02",X"E6",X"EA",X"02",X"EC",X"D3",X"D3",X"D3",
		X"EE",X"02",X"DE",X"E4",X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"EA",X"02",X"DC",X"FC",
		X"DA",X"02",X"DE",X"E4",X"02",X"E7",X"E9",X"EB",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"FC",X"FC",
		X"DA",X"02",X"E7",X"EB",X"02",X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DE",X"E4",X"02",X"DC",X"FC",
		X"DA",X"02",X"DE",X"E4",X"06",X"DE",X"E4",X"02",X"F0",X"FC",X"FC",X"FC",X"DA",X"05",X"DE",X"E4",
		X"05",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"E8",X"F4",
		X"E4",X"02",X"CE",X"FC",X"FC",X"FC",X"DA",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"E6",X"E8",
		X"E8",X"F4",X"E4",X"02",X"DC",X"00",X"62",X"02",X"01",X"13",X"01",X"01",X"01",X"02",X"01",X"04",
		X"03",X"13",X"06",X"04",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"06",X"04",X"03",X"10",X"03",X"06",X"04",X"03",
		X"10",X"03",X"06",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0C",X"03",X"01",X"01",X"01",
		X"01",X"01",X"01",X"07",X"04",X"0C",X"03",X"06",X"07",X"04",X"0C",X"03",X"06",X"04",X"01",X"01",
		X"01",X"04",X"0C",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"04",X"03",X"04",X"0F",X"03",X"03",
		X"04",X"03",X"04",X"0F",X"03",X"03",X"04",X"03",X"01",X"01",X"01",X"01",X"0F",X"01",X"01",X"01",
		X"03",X"04",X"03",X"19",X"04",X"03",X"19",X"04",X"03",X"01",X"01",X"01",X"01",X"0F",X"01",X"01",
		X"01",X"03",X"04",X"03",X"04",X"0F",X"03",X"03",X"04",X"03",X"04",X"0F",X"03",X"03",X"04",X"01",
		X"01",X"01",X"04",X"0C",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"07",X"04",X"0C",X"03",X"06",
		X"07",X"04",X"0C",X"03",X"06",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0C",X"03",X"01",
		X"01",X"01",X"01",X"01",X"01",X"04",X"03",X"10",X"03",X"06",X"04",X"03",X"10",X"03",X"06",X"04",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"06",X"04",X"03",X"13",X"06",X"04",X"02",X"01",X"13",X"01",X"01",X"01",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"1D",X"22",X"1D",X"39",X"40",X"20",X"40",X"3B",
		X"63",X"40",X"7C",X"40",X"83",X"43",X"9C",X"43",X"63",X"40",X"7C",X"40",X"63",X"43",X"7C",X"43",
		X"49",X"09",X"17",X"09",X"17",X"09",X"0E",X"E0",X"E0",X"E0",X"29",X"09",X"17",X"09",X"17",X"09",
		X"00",X"00",X"76",X"8A",X"13",X"94",X"0C",X"7B",X"8A",X"22",X"94",X"F4",X"84",X"8A",X"27",X"4C",
		X"F4",X"8E",X"8A",X"1C",X"4C",X"0C",X"80",X"AA",X"AA",X"BF",X"AA",X"80",X"0A",X"54",X"55",X"55",
		X"55",X"FF",X"5F",X"55",X"EA",X"FF",X"57",X"55",X"F5",X"57",X"FF",X"15",X"40",X"55",X"EA",X"AF",
		X"02",X"EA",X"FF",X"FF",X"AA",X"A7",X"8A",X"14",X"00",X"00",X"AC",X"8A",X"17",X"00",X"00",X"B2",
		X"8A",X"1A",X"00",X"00",X"B9",X"8A",X"1D",X"55",X"40",X"55",X"55",X"BF",X"AA",X"80",X"AA",X"AA",
		X"BF",X"AA",X"AA",X"80",X"AA",X"02",X"80",X"AA",X"AA",X"55",X"00",X"00",X"00",X"55",X"55",X"FD",
		X"AA",X"40",X"FC",X"DA",X"02",X"DE",X"D8",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D6",X"D8",
		X"D2",X"D2",X"D2",X"D2",X"D4",X"FC",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"D8",X"D2",X"D2",X"D2",
		X"D2",X"D4",X"FC",X"DA",X"02",X"DE",X"E4",X"08",X"DE",X"E4",X"05",X"DC",X"FC",X"FC",X"FC",X"FC",
		X"DA",X"02",X"DE",X"E4",X"05",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"E8",
		X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"EA",X"02",X"E7",X"D2",X"D2",X"D2",X"D2",X"EB",X"02",X"E7",
		X"EB",X"02",X"E6",X"EA",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"DE",X"F3",X"E9",X"E9",
		X"EB",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"0C",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"DE",
		X"E4",X"02",X"DE",X"E4",X"05",X"DE",X"E4",X"02",X"DE",X"F2",X"E8",X"E8",X"E8",X"EA",X"02",X"E6",
		X"EA",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"E7",X"EB",X"02",X"DE",
		X"E4",X"02",X"E6",X"EA",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"E9",X"EB",X"02",X"DE",
		X"E4",X"02",X"E7",X"E9",X"E9",X"E9",X"EB",X"02",X"DC",X"FC",X"DA",X"05",X"DE",X"E4",X"02",X"DE",
		X"E4",X"0C",X"DE",X"E4",X"08",X"DC",X"FC",X"FA",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"DE",
		X"F2",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"E6",X"E8",X"E8",X"EA",X"02",X"DE",X"F2",X"E8",X"E8",
		X"EA",X"02",X"E6",X"EA",X"02",X"DC",X"FC",X"FB",X"E9",X"E9",X"EB",X"02",X"E7",X"EB",X"02",X"E7",
		X"E9",X"E9",X"E9",X"E9",X"E9",X"EB",X"02",X"E7",X"E9",X"F5",X"E4",X"02",X"DE",X"F3",X"E9",X"E9",
		X"EB",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"12",X"DE",X"E4",X"02",X"DE",X"E4",X"05",X"DE",
		X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"E6",X"EA",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",
		X"EC",X"D3",X"D3",X"D3",X"EE",X"02",X"E7",X"EB",X"02",X"E7",X"EB",X"02",X"E6",X"EA",X"02",X"DE",
		X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E7",X"E9",X"E9",X"E9",X"F5",X"E4",X"02",
		X"DC",X"FC",X"FC",X"FC",X"DA",X"08",X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"DA",X"02",
		X"DE",X"E4",X"06",X"DE",X"E4",X"02",X"F0",X"FC",X"FC",X"FC",X"DA",X"02",X"E6",X"E8",X"E8",X"E8",
		X"EA",X"02",X"DE",X"E4",X"05",X"DC",X"FC",X"DA",X"02",X"DE",X"F2",X"E8",X"E8",X"E8",X"EA",X"02",
		X"DE",X"E4",X"02",X"CE",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"C0",X"C0",X"C0",X"E4",X"02",X"DE",
		X"F2",X"E8",X"E8",X"EA",X"02",X"DC",X"00",X"00",X"00",X"00",X"66",X"01",X"01",X"01",X"01",X"01",
		X"03",X"01",X"01",X"01",X"0B",X"01",X"01",X"07",X"06",X"03",X"03",X"0A",X"03",X"07",X"06",X"03",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"07",X"03",X"01",X"01",
		X"01",X"03",X"07",X"03",X"06",X"07",X"03",X"03",X"03",X"07",X"03",X"06",X"07",X"03",X"03",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",
		X"07",X"03",X"0D",X"06",X"03",X"07",X"03",X"0D",X"06",X"03",X"04",X"01",X"01",X"01",X"01",X"01",
		X"01",X"0D",X"03",X"01",X"01",X"01",X"03",X"04",X"03",X"10",X"03",X"03",X"03",X"04",X"03",X"10",
		X"01",X"01",X"01",X"03",X"03",X"04",X"03",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"04",
		X"07",X"15",X"04",X"07",X"15",X"04",X"03",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"04",
		X"03",X"10",X"01",X"01",X"01",X"03",X"03",X"04",X"03",X"10",X"03",X"03",X"03",X"04",X"01",X"01",
		X"01",X"01",X"01",X"01",X"0D",X"03",X"01",X"01",X"01",X"03",X"07",X"03",X"0D",X"06",X"03",X"07",
		X"03",X"0D",X"06",X"03",X"07",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"07",X"03",X"03",X"03",X"07",X"03",X"06",X"07",
		X"03",X"01",X"01",X"01",X"03",X"07",X"03",X"06",X"07",X"06",X"03",X"03",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"07",X"06",X"03",X"03",X"0A",X"03",X"08",X"01",X"01",
		X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"0B",X"01",X"01",X"F4",X"1D",X"22",X"1D",X"39",X"40",
		X"20",X"40",X"3B",X"65",X"40",X"7B",X"40",X"85",X"43",X"9B",X"43",X"65",X"40",X"7B",X"40",X"65",
		X"43",X"7B",X"43",X"42",X"16",X"0A",X"16",X"0A",X"16",X"0A",X"20",X"20",X"20",X"DE",X"E0",X"22",
		X"20",X"20",X"20",X"20",X"16",X"0A",X"16",X"0A",X"16",X"00",X"00",X"6F",X"8D",X"13",X"C4",X"0C",
		X"74",X"8D",X"1E",X"C4",X"F4",X"7C",X"8D",X"26",X"14",X"F4",X"86",X"8D",X"1D",X"14",X"0C",X"02",
		X"AA",X"AA",X"80",X"2A",X"02",X"40",X"55",X"7F",X"55",X"15",X"50",X"05",X"EA",X"FF",X"57",X"55",
		X"F5",X"FF",X"57",X"7F",X"55",X"05",X"EA",X"FF",X"FF",X"FF",X"EA",X"AF",X"AA",X"02",X"A2",X"8D",
		X"12",X"00",X"00",X"A7",X"8D",X"1D",X"00",X"00",X"AF",X"8D",X"21",X"00",X"00",X"B8",X"8D",X"2C",
		X"00",X"00",X"55",X"7F",X"55",X"D5",X"FF",X"AA",X"BF",X"AA",X"2A",X"A0",X"EA",X"FF",X"FF",X"AA",
		X"2A",X"A0",X"02",X"00",X"00",X"A0",X"AA",X"02",X"55",X"15",X"A0",X"2A",X"00",X"54",X"05",X"00",
		X"00",X"55",X"FD",X"40",X"FC",X"D0",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D6",X"E4",X"02",X"E7",
		X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D6",X"D8",X"D2",X"D2",X"D2",X"D2",
		X"D2",X"D2",X"D2",X"D4",X"FC",X"DA",X"07",X"DE",X"E4",X"0D",X"DE",X"E4",X"08",X"DC",X"FC",X"DA",
		X"02",X"E6",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"EA",X"02",X"E6",X"E8",
		X"E8",X"E8",X"EA",X"02",X"E7",X"EB",X"02",X"E6",X"EA",X"02",X"E6",X"EA",X"02",X"DC",X"FC",X"DA",
		X"02",X"DE",X"F3",X"E9",X"EB",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"F5",X"E4",X"02",X"E7",X"E9",
		X"E9",X"F5",X"E4",X"05",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",
		X"09",X"DE",X"E4",X"05",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"DE",X"E4",X"02",
		X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"E7",X"EB",
		X"02",X"E6",X"EA",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"EB",X"02",X"E7",X"EB",X"02",
		X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E7",X"E9",X"E9",X"E9",X"F5",X"E4",X"05",X"DE",X"E4",
		X"0E",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"06",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",
		X"02",X"E6",X"E8",X"E8",X"E8",X"EA",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"E8",X"F4",X"FC",X"DA",
		X"02",X"E7",X"EB",X"02",X"E6",X"E8",X"EA",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"EB",
		X"02",X"DE",X"F3",X"E9",X"E9",X"EB",X"02",X"DE",X"F3",X"E9",X"E9",X"E9",X"E9",X"F5",X"FC",X"DA",
		X"05",X"DE",X"C0",X"E4",X"0B",X"DE",X"E4",X"05",X"DE",X"E4",X"05",X"DC",X"FC",X"FA",X"E8",X"E8",
		X"EA",X"02",X"DE",X"C0",X"E4",X"02",X"E6",X"EA",X"02",X"EC",X"D3",X"D3",X"D3",X"EE",X"02",X"DE",
		X"E4",X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"EA",X"02",X"DC",X"FC",X"FB",X"E9",X"E9",
		X"EB",X"02",X"E7",X"E9",X"EB",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"E7",
		X"EB",X"02",X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"09",X"DE",
		X"E4",X"02",X"F0",X"FC",X"FC",X"FC",X"DA",X"05",X"DE",X"E4",X"05",X"DE",X"E4",X"02",X"DC",X"FC",
		X"DA",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"CE",X"FC",X"FC",X"FC",
		X"DA",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"DC",X"00",
		X"00",X"00",X"00",X"62",X"01",X"02",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"04",X"01",X"01",X"01",X"01",X"01",X"04",X"05",X"03",X"0B",X"03",X"03",
		X"03",X"04",X"05",X"03",X"0B",X"01",X"01",X"01",X"03",X"03",X"04",X"03",X"01",X"01",X"01",X"01",
		X"01",X"0B",X"06",X"03",X"04",X"03",X"10",X"06",X"03",X"04",X"03",X"10",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"04",X"03",X"01",X"01",X"01",X"01",X"0F",X"0A",X"03",X"04",X"0F",
		X"0A",X"01",X"01",X"01",X"04",X"0C",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"07",X"04",X"0C",
		X"03",X"03",X"03",X"07",X"04",X"0C",X"03",X"03",X"03",X"04",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"0C",X"03",X"01",X"01",X"01",X"03",X"04",X"07",X"15",X"04",X"07",X"15",X"04",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"0C",X"03",X"01",X"01",X"01",X"03",X"07",X"04",X"0C",X"03",X"03",
		X"03",X"07",X"04",X"0C",X"03",X"03",X"03",X"04",X"01",X"01",X"01",X"04",X"0C",X"01",X"01",X"01",
		X"03",X"01",X"01",X"01",X"04",X"03",X"04",X"0F",X"0A",X"03",X"01",X"01",X"01",X"01",X"0F",X"0A",
		X"03",X"10",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"03",X"10",X"06",X"03",
		X"04",X"03",X"01",X"01",X"01",X"01",X"01",X"0B",X"06",X"03",X"04",X"05",X"03",X"0B",X"01",X"01",
		X"01",X"03",X"03",X"04",X"05",X"03",X"0B",X"03",X"03",X"03",X"04",X"01",X"02",X"01",X"01",X"03",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"01",X"01",X"01",X"01",
		X"01",X"00",X"00",X"00",X"F2",X"40",X"2D",X"1D",X"22",X"1D",X"39",X"40",X"20",X"64",X"40",X"78",
		X"40",X"84",X"43",X"98",X"43",X"64",X"40",X"78",X"40",X"64",X"43",X"78",X"43",X"51",X"90",X"15",
		X"54",X"0C",X"57",X"90",X"1E",X"54",X"F4",X"57",X"90",X"1E",X"54",X"F4",X"5F",X"90",X"15",X"54",
		X"0C",X"EA",X"FF",X"AB",X"FA",X"AA",X"AA",X"EA",X"FF",X"57",X"55",X"55",X"D5",X"57",X"55",X"AA",
		X"AA",X"BF",X"FA",X"BF",X"AA",X"79",X"90",X"22",X"00",X"00",X"82",X"90",X"25",X"00",X"00",X"82",
		X"90",X"25",X"00",X"00",X"92",X"90",X"28",X"00",X"00",X"05",X"00",X"00",X"54",X"05",X"54",X"7F",
		X"F5",X"0B",X"0A",X"00",X"00",X"A8",X"0A",X"A8",X"BF",X"FA",X"AB",X"AA",X"AA",X"82",X"AA",X"00",
		X"A0",X"AA",X"55",X"41",X"55",X"00",X"A0",X"02",X"40",X"F5",X"57",X"BF",X"40",X"FC",X"D0",X"D2",
		X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D4",X"FC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"DC",
		X"FC",X"FC",X"FC",X"FC",X"D0",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D4",X"FC",X"DA",X"09",
		X"DC",X"FC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"FC",X"FC",X"FC",X"DA",X"08",X"DC",
		X"FC",X"DA",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"E7",X"D2",X"D2",X"EB",X"02",X"DE",
		X"E4",X"02",X"E7",X"D2",X"D2",X"D2",X"D2",X"EB",X"02",X"E6",X"E8",X"E8",X"E8",X"EA",X"02",X"DC",
		X"FC",X"DA",X"02",X"E7",X"E9",X"E9",X"E9",X"F5",X"E4",X"07",X"DE",X"E4",X"09",X"DE",X"F3",X"E9",
		X"E9",X"EB",X"02",X"DC",X"FC",X"DA",X"06",X"DE",X"E4",X"02",X"E6",X"EA",X"02",X"E6",X"E8",X"F4",
		X"F2",X"E8",X"EA",X"02",X"E6",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"05",X"DC",X"FC",X"DA",X"02",
		X"E6",X"E8",X"EA",X"02",X"E7",X"EB",X"02",X"DE",X"E4",X"02",X"E7",X"E9",X"E9",X"E9",X"E9",X"EB",
		X"02",X"E7",X"E9",X"F5",X"E4",X"02",X"E7",X"EB",X"02",X"E6",X"EA",X"02",X"DC",X"FC",X"DA",X"02",
		X"DE",X"C0",X"E4",X"05",X"DE",X"E4",X"0B",X"DE",X"E4",X"05",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",
		X"02",X"DE",X"C0",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"F2",X"E8",X"E8",X"EA",X"02",X"E6",X"E8",
		X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"DC",X"FC",X"DA",
		X"02",X"E7",X"E9",X"EB",X"02",X"E7",X"E9",X"E9",X"F5",X"F3",X"E9",X"E9",X"EB",X"02",X"E7",X"E9",
		X"E9",X"F5",X"E4",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"F5",X"E4",X"02",X"DC",X"FC",X"DA",
		X"09",X"DE",X"E4",X"08",X"DE",X"E4",X"08",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"E6",X"E8",
		X"E8",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"EC",X"D3",X"D3",X"D3",X"EE",X"02",X"DE",X"E4",
		X"02",X"E6",X"E8",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"F3",
		X"E9",X"E9",X"E9",X"EB",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"E7",X"EB",
		X"02",X"E7",X"E9",X"E9",X"F5",X"E4",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",
		X"09",X"F0",X"FC",X"FC",X"FC",X"DA",X"08",X"DE",X"E4",X"05",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",
		X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"CE",X"FC",X"FC",X"FC",X"DA",X"02",X"E6",X"E8",
		X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"00",X"00",X"00",X"00",X"62",
		X"01",X"02",X"01",X"01",X"01",X"01",X"0F",X"01",X"01",X"01",X"02",X"01",X"04",X"07",X"0F",X"06",
		X"04",X"07",X"01",X"01",X"01",X"07",X"01",X"01",X"01",X"01",X"01",X"06",X"04",X"01",X"01",X"01",
		X"01",X"03",X"03",X"07",X"05",X"03",X"01",X"01",X"01",X"04",X"04",X"03",X"03",X"07",X"05",X"03",
		X"03",X"04",X"04",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"03",X"01",X"01",X"01",X"03",X"04",X"04",X"0F",X"03",X"06",X"04",X"04",X"0F",X"03",X"06",X"04",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0C",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"04",
		X"07",X"12",X"03",X"04",X"07",X"12",X"03",X"04",X"03",X"01",X"01",X"01",X"01",X"12",X"01",X"01",
		X"01",X"04",X"03",X"16",X"07",X"03",X"16",X"07",X"03",X"01",X"01",X"01",X"01",X"12",X"01",X"01",
		X"01",X"04",X"07",X"12",X"03",X"04",X"07",X"12",X"03",X"04",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"0C",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"04",X"04",X"0F",X"03",X"06",X"04",X"04",
		X"0F",X"03",X"06",X"04",X"04",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"04",X"04",X"03",X"03",X"07",X"05",X"03",X"03",X"04",
		X"01",X"01",X"01",X"01",X"03",X"03",X"07",X"05",X"03",X"01",X"01",X"01",X"04",X"07",X"01",X"01",
		X"01",X"07",X"01",X"01",X"01",X"01",X"01",X"06",X"04",X"07",X"0F",X"06",X"04",X"01",X"02",X"01",
		X"01",X"01",X"01",X"0F",X"01",X"01",X"01",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"EF",X"1C",X"36",
		X"EF",X"20",X"15",X"EF",X"21",X"13",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",X"EF",X"1C",
		X"36",X"EF",X"20",X"16",X"EF",X"21",X"14",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",X"EF",
		X"1C",X"36",X"EF",X"20",X"17",X"EF",X"21",X"15",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",
		X"EF",X"1C",X"36",X"EF",X"20",X"18",X"EF",X"21",X"16",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",
		X"F5",X"EF",X"1C",X"36",X"EF",X"20",X"18",X"EF",X"21",X"17",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",
		X"C9",X"F5",X"EF",X"1C",X"36",X"EF",X"20",X"19",X"EF",X"21",X"18",X"21",X"BC",X"4E",X"CB",X"DE",
		X"F1",X"C9",X"F5",X"EF",X"1C",X"36",X"EF",X"20",X"1A",X"EF",X"21",X"19",X"21",X"BC",X"4E",X"CB",
		X"DE",X"F1",X"C9",X"EE",X"64",X"40",X"7C",X"40",X"84",X"43",X"9C",X"43",X"64",X"40",X"7C",X"40",
		X"64",X"43",X"7C",X"43",X"1D",X"22",X"40",X"20",X"1D",X"39",X"40",X"3B",X"C0",X"93",X"14",X"8C",
		X"0C",X"C5",X"93",X"1D",X"8C",X"F4",X"CE",X"93",X"2A",X"74",X"F4",X"D9",X"93",X"15",X"74",X"0C",
		X"80",X"AA",X"BE",X"FA",X"AA",X"00",X"00",X"50",X"FD",X"55",X"F5",X"D5",X"57",X"55",X"EA",X"FF",
		X"57",X"D5",X"5F",X"FD",X"15",X"50",X"01",X"50",X"55",X"EA",X"AF",X"FE",X"2A",X"A8",X"AA",X"F3",
		X"93",X"15",X"00",X"00",X"F9",X"93",X"18",X"00",X"00",X"FF",X"93",X"19",X"00",X"00",X"06",X"94",
		X"1C",X"00",X"00",X"55",X"50",X"41",X"55",X"FD",X"AA",X"AA",X"A0",X"82",X"AA",X"FE",X"AA",X"AA",
		X"AF",X"02",X"2A",X"A0",X"AA",X"AA",X"55",X"5F",X"01",X"00",X"50",X"55",X"BF",X"3A",X"70",X"4C",
		X"FE",X"02",X"20",X"07",X"3A",X"13",X"4E",X"FE",X"08",X"30",X"05",X"21",X"2A",X"94",X"18",X"03",
		X"21",X"32",X"94",X"CD",X"A1",X"94",X"21",X"00",X"40",X"C9",X"CC",X"87",X"C1",X"8A",X"C3",X"8D",
		X"9C",X"90",X"5F",X"99",X"D2",X"9B",X"43",X"9E",X"AE",X"A0",X"21",X"68",X"22",X"18",X"03",X"21",
		X"90",X"22",X"E5",X"3A",X"70",X"4C",X"FE",X"02",X"20",X"07",X"3A",X"13",X"4E",X"FE",X"08",X"30",
		X"05",X"21",X"6A",X"94",X"18",X"03",X"21",X"72",X"94",X"CD",X"A1",X"94",X"FD",X"21",X"00",X"00",
		X"FD",X"09",X"21",X"00",X"40",X"DD",X"21",X"16",X"4E",X"C9",X"46",X"89",X"3A",X"8C",X"33",X"8F",
		X"0F",X"92",X"E1",X"9A",X"4B",X"9D",X"B7",X"9F",X"21",X"A2",X"C5",X"21",X"99",X"94",X"CD",X"A1",
		X"94",X"0A",X"47",X"3A",X"0E",X"4E",X"B8",X"C1",X"DA",X"8E",X"94",X"C3",X"42",X"0B",X"3A",X"FD",
		X"4D",X"FE",X"05",X"DA",X"48",X"0B",X"C3",X"42",X"0B",X"37",X"8A",X"2A",X"8D",X"24",X"90",X"93",
		X"93",X"3A",X"13",X"4E",X"E5",X"FE",X"0D",X"F2",X"B8",X"94",X"21",X"C3",X"94",X"D7",X"E1",X"87",
		X"4F",X"06",X"00",X"09",X"4E",X"23",X"46",X"C9",X"D6",X"0D",X"D6",X"08",X"F2",X"BA",X"94",X"C6",
		X"0D",X"18",X"E7",X"00",X"00",X"01",X"01",X"02",X"02",X"03",X"03",X"00",X"01",X"02",X"03",X"00",
		X"01",X"02",X"03",X"03",X"03",X"02",X"01",X"3A",X"70",X"4C",X"FE",X"03",X"CC",X"90",X"B3",X"21",
		X"2D",X"95",X"CD",X"A1",X"94",X"11",X"34",X"4E",X"69",X"60",X"4E",X"23",X"46",X"23",X"1A",X"FE",
		X"14",X"28",X"04",X"FE",X"40",X"20",X"08",X"02",X"13",X"3E",X"03",X"A3",X"20",X"EC",X"C9",X"3E",
		X"40",X"12",X"02",X"18",X"F3",X"3A",X"70",X"4C",X"FE",X"03",X"CC",X"90",X"B3",X"21",X"2D",X"95",
		X"CD",X"A1",X"94",X"11",X"34",X"4E",X"69",X"60",X"4E",X"23",X"46",X"23",X"0A",X"FE",X"14",X"28",
		X"04",X"FE",X"40",X"20",X"01",X"12",X"13",X"3E",X"03",X"A3",X"20",X"EC",X"C9",X"40",X"8A",X"33",
		X"8D",X"2D",X"90",X"94",X"93",X"48",X"8A",X"3B",X"8D",X"35",X"90",X"9C",X"93",X"C5",X"D5",X"21",
		X"2D",X"95",X"CD",X"A1",X"94",X"60",X"69",X"5E",X"23",X"56",X"EB",X"CB",X"D4",X"3A",X"7E",X"44",
		X"BE",X"20",X"02",X"3E",X"00",X"77",X"EB",X"23",X"5E",X"23",X"56",X"CB",X"D2",X"12",X"23",X"5E",
		X"23",X"56",X"CB",X"D2",X"12",X"23",X"5E",X"23",X"56",X"CB",X"D2",X"12",X"D1",X"C1",X"3E",X"10",
		X"BE",X"C9",X"3A",X"2E",X"4D",X"18",X"03",X"3A",X"2F",X"4D",X"F5",X"C5",X"E5",X"21",X"91",X"95",
		X"CD",X"A1",X"94",X"69",X"60",X"ED",X"5F",X"E6",X"06",X"D7",X"5F",X"23",X"56",X"E1",X"C1",X"F1",
		X"C9",X"38",X"8A",X"2B",X"8D",X"25",X"90",X"A4",X"93",X"CA",X"CD",X"22",X"3A",X"02",X"4E",X"A7",
		X"28",X"07",X"FE",X"10",X"3E",X"01",X"C2",X"CD",X"22",X"3A",X"13",X"4E",X"FE",X"15",X"F2",X"BC",
		X"95",X"4F",X"06",X"00",X"21",X"C7",X"95",X"09",X"7E",X"C3",X"CD",X"22",X"D6",X"15",X"D6",X"10",
		X"F2",X"BE",X"95",X"C6",X"15",X"18",X"EA",X"07",X"16",X"1D",X"07",X"14",X"09",X"07",X"14",X"12",
		X"07",X"1D",X"14",X"16",X"18",X"1E",X"19",X"18",X"15",X"19",X"1D",X"12",X"07",X"16",X"1D",X"07",
		X"14",X"16",X"07",X"14",X"1D",X"07",X"1D",X"14",X"16",X"18",X"18",X"18",X"18",X"1D",X"1D",X"1D",
		X"1D",X"3A",X"13",X"4E",X"FE",X"03",X"F2",X"20",X"23",X"21",X"0D",X"96",X"CD",X"A1",X"94",X"21",
		X"00",X"44",X"0A",X"03",X"A7",X"CA",X"20",X"23",X"D7",X"CB",X"F6",X"18",X"F5",X"50",X"8A",X"43",
		X"8D",X"50",X"8A",X"43",X"8D",X"78",X"FE",X"0A",X"CC",X"3A",X"96",X"FE",X"0B",X"CC",X"28",X"96",
		X"FE",X"06",X"CC",X"FE",X"96",X"C3",X"DF",X"2A",X"C5",X"E5",X"E1",X"C1",X"3A",X"80",X"50",X"E6",
		X"30",X"FE",X"30",X"78",X"C0",X"3E",X"20",X"06",X"20",X"C9",X"C5",X"E5",X"21",X"45",X"96",X"CD",
		X"E9",X"96",X"E1",X"C1",X"C9",X"09",X"20",X"F5",X"41",X"09",X"21",X"15",X"42",X"09",X"22",X"F6",
		X"41",X"09",X"23",X"16",X"42",X"FF",X"3A",X"DA",X"4F",X"EF",X"64",X"96",X"65",X"96",X"86",X"96",
		X"A7",X"96",X"C8",X"96",X"C9",X"21",X"64",X"80",X"22",X"00",X"4D",X"21",X"2C",X"2E",X"22",X"0A",
		X"4D",X"22",X"31",X"4D",X"21",X"00",X"01",X"22",X"14",X"4D",X"22",X"1E",X"4D",X"3E",X"02",X"32",
		X"28",X"4D",X"32",X"2C",X"4D",X"C9",X"21",X"7C",X"80",X"22",X"02",X"4D",X"21",X"2F",X"2E",X"22",
		X"0C",X"4D",X"22",X"33",X"4D",X"21",X"01",X"00",X"22",X"16",X"4D",X"22",X"20",X"4D",X"3E",X"01",
		X"32",X"29",X"4D",X"32",X"2D",X"4D",X"C9",X"21",X"7C",X"90",X"22",X"04",X"4D",X"21",X"2F",X"30",
		X"22",X"0E",X"4D",X"22",X"35",X"4D",X"21",X"FF",X"00",X"22",X"18",X"4D",X"22",X"22",X"4D",X"3E",
		X"03",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"C9",X"21",X"7C",X"70",X"22",X"06",X"4D",X"21",X"2F",
		X"2C",X"22",X"10",X"4D",X"22",X"37",X"4D",X"21",X"FF",X"00",X"22",X"1A",X"4D",X"22",X"24",X"4D",
		X"3E",X"03",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"C9",X"7E",X"FE",X"FF",X"28",X"0F",X"47",X"23",
		X"7E",X"23",X"5E",X"23",X"56",X"12",X"78",X"CB",X"D2",X"12",X"23",X"18",X"EC",X"C9",X"3E",X"00",
		X"32",X"00",X"4F",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"34",X"3E",X"CD",
		X"49",X"97",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",
		X"E5",X"FD",X"E5",X"CD",X"4C",X"3E",X"CD",X"17",X"3F",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",
		X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"01",X"80",X"CD",X"8F",X"06",
		X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"3A",X"01",X"4F",X"3C",X"E6",X"1F",X"32",
		X"01",X"4F",X"E6",X"07",X"4F",X"CB",X"81",X"06",X"00",X"DD",X"21",X"D9",X"98",X"CB",X"47",X"CA",
		X"E7",X"97",X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"36",X"87",X"DD",X"6E",X"08",X"DD",
		X"66",X"09",X"36",X"87",X"DD",X"6E",X"10",X"DD",X"66",X"11",X"36",X"87",X"DD",X"6E",X"18",X"DD",
		X"66",X"19",X"36",X"87",X"DD",X"6E",X"20",X"DD",X"66",X"21",X"36",X"87",X"DD",X"6E",X"28",X"DD",
		X"66",X"29",X"3E",X"67",X"BD",X"20",X"04",X"36",X"8A",X"18",X"02",X"36",X"87",X"DD",X"6E",X"30",
		X"DD",X"66",X"31",X"36",X"8A",X"DD",X"6E",X"38",X"DD",X"66",X"39",X"36",X"81",X"DD",X"6E",X"40",
		X"DD",X"66",X"41",X"36",X"81",X"DD",X"6E",X"48",X"DD",X"66",X"49",X"36",X"81",X"DD",X"6E",X"50",
		X"DD",X"66",X"51",X"36",X"81",X"DD",X"6E",X"58",X"DD",X"66",X"59",X"36",X"81",X"DD",X"6E",X"60",
		X"DD",X"66",X"61",X"3E",X"63",X"BD",X"20",X"04",X"36",X"84",X"18",X"02",X"36",X"81",X"DD",X"6E",
		X"68",X"DD",X"66",X"69",X"36",X"84",X"C9",X"0D",X"AF",X"B9",X"FA",X"EF",X"97",X"06",X"FF",X"0D",
		X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"35",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"36",
		X"88",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"35",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"36",X"88",
		X"DD",X"6E",X"10",X"DD",X"66",X"11",X"35",X"DD",X"6E",X"12",X"DD",X"66",X"13",X"36",X"88",X"DD",
		X"6E",X"18",X"DD",X"66",X"19",X"35",X"DD",X"6E",X"1A",X"DD",X"66",X"1B",X"36",X"88",X"DD",X"6E",
		X"20",X"DD",X"66",X"21",X"35",X"DD",X"6E",X"22",X"DD",X"66",X"23",X"36",X"88",X"DD",X"6E",X"28",
		X"DD",X"66",X"29",X"35",X"DD",X"6E",X"2A",X"DD",X"66",X"2B",X"3E",X"67",X"BD",X"20",X"04",X"36",
		X"8B",X"18",X"02",X"36",X"88",X"DD",X"6E",X"30",X"DD",X"66",X"31",X"35",X"DD",X"6E",X"32",X"DD",
		X"66",X"33",X"36",X"8B",X"DD",X"6E",X"38",X"DD",X"66",X"39",X"35",X"DD",X"6E",X"3A",X"DD",X"66",
		X"3B",X"36",X"82",X"DD",X"6E",X"40",X"DD",X"66",X"41",X"35",X"DD",X"6E",X"42",X"DD",X"66",X"43",
		X"36",X"82",X"DD",X"6E",X"48",X"DD",X"66",X"49",X"35",X"DD",X"6E",X"4A",X"DD",X"66",X"4B",X"36",
		X"82",X"DD",X"6E",X"50",X"DD",X"66",X"51",X"35",X"DD",X"6E",X"52",X"DD",X"66",X"53",X"36",X"82",
		X"DD",X"6E",X"58",X"DD",X"66",X"59",X"35",X"DD",X"6E",X"5A",X"DD",X"66",X"5B",X"36",X"82",X"DD",
		X"6E",X"60",X"DD",X"66",X"61",X"35",X"DD",X"6E",X"62",X"DD",X"66",X"63",X"3E",X"63",X"BD",X"20",
		X"04",X"36",X"83",X"18",X"02",X"36",X"82",X"DD",X"6E",X"68",X"DD",X"66",X"69",X"35",X"DD",X"6E",
		X"6A",X"DD",X"66",X"6B",X"36",X"83",X"C9",X"67",X"43",X"47",X"43",X"27",X"43",X"07",X"43",X"E7",
		X"42",X"C7",X"42",X"A7",X"42",X"87",X"42",X"67",X"42",X"47",X"42",X"27",X"42",X"07",X"42",X"E7",
		X"41",X"C7",X"41",X"A7",X"41",X"87",X"41",X"67",X"41",X"47",X"41",X"27",X"41",X"07",X"41",X"E7",
		X"40",X"C7",X"40",X"A7",X"40",X"87",X"40",X"67",X"40",X"66",X"40",X"65",X"40",X"64",X"40",X"63",
		X"40",X"83",X"40",X"A3",X"40",X"C3",X"40",X"E3",X"40",X"03",X"41",X"23",X"41",X"43",X"41",X"63",
		X"41",X"83",X"41",X"A3",X"41",X"C3",X"41",X"E3",X"41",X"03",X"42",X"23",X"42",X"43",X"42",X"63",
		X"42",X"83",X"42",X"A3",X"42",X"C3",X"42",X"E3",X"42",X"03",X"43",X"23",X"43",X"43",X"43",X"63",
		X"43",X"64",X"43",X"65",X"43",X"66",X"43",X"67",X"43",X"64",X"43",X"65",X"43",X"66",X"43",X"67",
		X"43",X"64",X"43",X"65",X"43",X"66",X"43",X"67",X"43",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"FC",X"D0",X"EF",X"02",X"ED",X"D2",X"D2",X"EF",X"02",X"ED",X"D4",X"FC",X"FC",X"FC",X"DA",X"02",
		X"DC",X"FC",X"FC",X"FC",X"D0",X"EF",X"02",X"ED",X"D2",X"D6",X"E4",X"02",X"ED",X"D2",X"D2",X"D4",
		X"02",X"DA",X"09",X"F7",X"D2",X"D2",X"D2",X"EB",X"02",X"F7",X"D2",X"D2",X"D2",X"EB",X"05",X"DE",
		X"E4",X"05",X"DC",X"02",X"DA",X"02",X"E6",X"E8",X"EA",X"02",X"E6",X"EA",X"0E",X"E6",X"EA",X"02",
		X"E7",X"EB",X"02",X"E6",X"EA",X"02",X"DC",X"02",X"DA",X"02",X"DE",X"FC",X"E4",X"02",X"DE",X"E4",
		X"02",X"F6",X"D3",X"D3",X"D3",X"EA",X"02",X"F6",X"D3",X"D3",X"D3",X"EA",X"02",X"DE",X"E4",X"05",
		X"DE",X"E4",X"02",X"DC",X"02",X"DA",X"02",X"DE",X"FC",X"E4",X"02",X"DE",X"E4",X"02",X"DC",X"FC",
		X"FC",X"FC",X"DA",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"F2",X"E8",X"E8",X"EA",X"02",
		X"E7",X"EB",X"02",X"DC",X"02",X"DA",X"02",X"E7",X"E9",X"EB",X"02",X"E7",X"EB",X"02",X"E7",X"D2",
		X"D2",X"D2",X"EB",X"02",X"E7",X"D2",X"D2",X"D2",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"EB",X"05",
		X"DC",X"02",X"DA",X"1B",X"E6",X"EA",X"02",X"DC",X"02",X"DA",X"02",X"E6",X"E8",X"F8",X"02",X"F6",
		X"E8",X"E8",X"E8",X"E8",X"F8",X"02",X"F6",X"E8",X"F8",X"02",X"F6",X"E8",X"EA",X"02",X"E6",X"F8",
		X"02",X"F6",X"E8",X"E8",X"F4",X"E4",X"02",X"DC",X"02",X"DA",X"02",X"DE",X"FC",X"E4",X"02",X"F7",
		X"E9",X"E9",X"F5",X"F3",X"F9",X"02",X"F7",X"E9",X"F9",X"02",X"F7",X"E9",X"EB",X"02",X"DE",X"E4",
		X"02",X"F7",X"E9",X"E9",X"F5",X"E4",X"02",X"DC",X"02",X"DA",X"02",X"DE",X"FC",X"E4",X"05",X"DE",
		X"E4",X"0B",X"DE",X"E4",X"05",X"DE",X"E4",X"02",X"DC",X"02",X"DA",X"02",X"DE",X"FC",X"E4",X"02",
		X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"EC",X"D3",X"D3",X"D3",X"EE",X"02",X"E6",X"EA",X"02",X"DE",
		X"E4",X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"DC",X"02",X"DA",X"02",X"E7",X"E9",X"EB",X"02",
		X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E7",
		X"EB",X"02",X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DC",X"02",X"DA",X"06",X"DE",X"E4",X"05",X"F0",
		X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"E4",X"05",X"DE",X"E4",X"05",X"DC",X"02",X"FA",X"E8",X"E8",
		X"EA",X"02",X"F6",X"F4",X"F2",X"E8",X"E8",X"EA",X"02",X"CE",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",
		X"F2",X"E8",X"E8",X"EA",X"02",X"DE",X"F2",X"EA",X"02",X"F6",X"E8",X"D5",X"00",X"00",X"00",X"00",
		X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"62",X"01",X"18",X"01",X"01",X"01",X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"04",
		X"03",X"0C",X"03",X"01",X"01",X"01",X"03",X"04",X"04",X"03",X"0C",X"06",X"03",X"04",X"04",X"03",
		X"0C",X"07",X"02",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"04",X"04",
		X"0F",X"03",X"06",X"04",X"04",X"0F",X"03",X"06",X"04",X"04",X"01",X"01",X"01",X"0C",X"03",X"01",
		X"01",X"01",X"03",X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"04",X"03",X"0C",X"03",X"03",
		X"03",X"04",X"01",X"01",X"01",X"01",X"03",X"0C",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"07",
		X"17",X"09",X"17",X"06",X"01",X"01",X"01",X"01",X"03",X"0C",X"01",X"01",X"01",X"03",X"01",X"01",
		X"01",X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",
		X"04",X"01",X"01",X"01",X"0C",X"03",X"01",X"01",X"01",X"03",X"04",X"04",X"0F",X"03",X"06",X"04",
		X"04",X"0F",X"03",X"06",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"04",
		X"04",X"03",X"0C",X"07",X"02",X"04",X"04",X"03",X"0C",X"06",X"03",X"04",X"04",X"03",X"0C",X"03",
		X"01",X"01",X"01",X"03",X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"01",X"18",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"FC",X"D0",X"D2",X"D2",X"D2",X"D2",X"D6",X"E4",X"02",X"DE",X"D8",X"D2",X"D2",
		X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D6",X"E4",X"02",X"DE",X"D8",X"D2",X"D2",X"D2",X"D2",X"D2",
		X"D2",X"D2",X"D4",X"FC",X"DA",X"05",X"DE",X"E4",X"02",X"DE",X"E4",X"09",X"DE",X"E4",X"02",X"DE",
		X"E4",X"08",X"DC",X"FC",X"DA",X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"E6",
		X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"E8",
		X"EA",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DE",
		X"C0",X"C0",X"C0",X"C0",X"E4",X"02",X"E7",X"EB",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",
		X"EB",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DE",
		X"C0",X"C0",X"C0",X"C0",X"E4",X"0E",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E7",X"EB",X"02",
		X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"E9",X"EB",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"E8",
		X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"0F",X"DE",X"F3",X"E9",
		X"E9",X"E9",X"E9",X"F5",X"F3",X"E9",X"E9",X"EB",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",
		X"E6",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"05",
		X"DE",X"E4",X"05",X"DC",X"FC",X"DA",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"F5",X"F3",
		X"E9",X"E9",X"E9",X"E9",X"E9",X"EB",X"02",X"DE",X"E4",X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",
		X"E6",X"EA",X"02",X"DC",X"FC",X"DA",X"09",X"DE",X"E4",X"08",X"DE",X"E4",X"02",X"DE",X"E4",X"02",
		X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"FA",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"EA",
		X"02",X"DE",X"E4",X"02",X"EC",X"D3",X"D3",X"D3",X"EE",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",
		X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"FB",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"EB",
		X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"E7",X"EB",X"02",X"DE",X"E4",X"02",
		X"E7",X"EB",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"DA",X"0C",X"DC",X"FC",X"FC",X"FC",X"DA",X"05",
		X"DE",X"E4",X"08",X"DC",X"FC",X"DA",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"EA",
		X"02",X"CE",X"FC",X"FC",X"FC",X"DA",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"E6",X"E8",X"E8",
		X"E8",X"E8",X"E8",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"01",X"01",X"07",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"06",X"01",X"01",X"02",X"01",X"01",X"04",X"03",X"06",X"07",
		X"06",X"06",X"04",X"03",X"06",X"07",X"06",X"06",X"04",X"03",X"06",X"07",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"03",X"06",X"07",X"0C",X"04",X"03",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0C",X"04",X"03",X"10",
		X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"04",X"03",X"10",X"03",X"03",X"03",X"04",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"0C",X"03",X"03",X"03",X"0B",X"0C",X"03",X"03",X"03",X"0B",X"0C",
		X"03",X"03",X"03",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"01",X"01",X"01",X"01",
		X"01",X"01",X"04",X"20",X"20",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"01",X"01",X"01",
		X"01",X"01",X"01",X"0B",X"0C",X"03",X"03",X"03",X"0B",X"0C",X"03",X"03",X"03",X"04",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"0C",X"03",X"03",X"03",X"04",X"03",X"10",X"03",X"03",X"03",X"04",
		X"03",X"10",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"04",X"03",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0C",X"04",X"03",X"06",X"07",X"0C",X"04",X"03",
		X"06",X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"03",
		X"06",X"07",X"06",X"06",X"04",X"03",X"06",X"07",X"06",X"06",X"04",X"01",X"01",X"07",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"06",X"01",X"01",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"FC",X"D0",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",
		X"D2",X"D6",X"D8",X"D2",X"D2",X"D2",X"D2",X"D2",X"EB",X"02",X"DE",X"D8",X"D2",X"D2",X"D2",X"D2",
		X"D2",X"D2",X"D2",X"D4",X"FC",X"DA",X"0C",X"DE",X"E4",X"08",X"DE",X"E4",X"08",X"DC",X"FC",X"DA",
		X"02",X"E6",X"EA",X"02",X"E6",X"EA",X"02",X"E6",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",
		X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"E8",X"EA",X"02",X"DC",X"FC",X"DA",
		X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DE",X"C0",X"E4",X"02",X"DE",X"E4",X"02",X"DE",X"C0",
		X"C0",X"C0",X"E4",X"02",X"DE",X"E4",X"02",X"E7",X"E9",X"E9",X"E9",X"EB",X"02",X"DC",X"FC",X"DA",
		X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DE",X"C0",X"E4",X"02",X"E7",X"EB",X"02",X"DE",X"C0",
		X"C0",X"C0",X"E4",X"02",X"DE",X"E4",X"08",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",
		X"02",X"E7",X"E9",X"EB",X"05",X"E7",X"E9",X"E9",X"E9",X"EB",X"02",X"DE",X"E4",X"02",X"E6",X"E8",
		X"E8",X"E8",X"EA",X"02",X"DC",X"FC",X"DA",X"02",X"E7",X"EB",X"02",X"E7",X"EB",X"06",X"E6",X"EA",
		X"08",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"EB",X"02",X"DC",X"FC",X"DA",X"08",X"E6",X"E8",
		X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"E8",X"EA",X"0B",X"DC",X"FC",X"DA",X"02",X"E6",
		X"EA",X"02",X"E6",X"EA",X"02",X"E7",X"E9",X"EB",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",
		X"EB",X"02",X"E6",X"E8",X"EA",X"02",X"E6",X"E8",X"E8",X"EA",X"02",X"DC",X"FC",X"DA",X"02",X"DE",
		X"E4",X"02",X"DE",X"E4",X"0F",X"E7",X"E9",X"EB",X"02",X"E7",X"E9",X"F5",X"E4",X"02",X"DC",X"FC",
		X"DA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"EA",X"02",X"EC",X"D3",X"D3",X"D3",
		X"EE",X"02",X"E6",X"EA",X"08",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"E7",X"EB",X"02",X"E7",
		X"EB",X"02",X"DE",X"C0",X"E4",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"E6",
		X"EA",X"02",X"E6",X"EA",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"DA",X"08",X"DE",X"C0",X"E4",X"02",
		X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"05",X"DC",
		X"FC",X"F2",X"E8",X"E8",X"E8",X"EA",X"02",X"E6",X"E8",X"F4",X"C0",X"E4",X"02",X"CE",X"FC",X"FC",
		X"FC",X"DA",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"01",X"01",X"01",X"01",X"01",X"04",X"03",
		X"03",X"04",X"03",X"06",X"03",X"06",X"04",X"03",X"03",X"04",X"03",X"06",X"03",X"06",X"04",X"03",
		X"03",X"04",X"03",X"06",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"03",X"03",X"04",X"01",
		X"01",X"01",X"06",X"03",X"06",X"04",X"03",X"03",X"0D",X"03",X"06",X"04",X"01",X"01",X"01",X"01",
		X"01",X"01",X"0D",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"03",X"03",X"11",
		X"05",X"04",X"03",X"03",X"11",X"05",X"04",X"03",X"03",X"11",X"01",X"01",X"03",X"04",X"03",X"03",
		X"13",X"03",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"08",X"20",X"1C",
		X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"04",X"03",X"03",X"13",X"03",X"04",
		X"03",X"03",X"11",X"01",X"01",X"03",X"04",X"03",X"03",X"11",X"05",X"04",X"03",X"03",X"11",X"05",
		X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"0D",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"04",X"03",X"03",X"0D",X"03",X"06",X"04",X"03",X"03",X"04",X"01",X"01",X"01",X"06",X"03",
		X"06",X"04",X"03",X"03",X"04",X"03",X"06",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"03",
		X"03",X"04",X"03",X"06",X"03",X"06",X"04",X"03",X"03",X"04",X"03",X"06",X"03",X"06",X"04",X"01",
		X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"04",
		X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"FC",
		X"D0",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"F5",X"C0",X"C0",X"C0",X"C0",X"E4",X"02",
		X"DE",X"C0",X"C0",X"C0",X"C0",X"C0",X"D8",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D4",X"FC",
		X"DA",X"09",X"DE",X"C0",X"C0",X"C0",X"C0",X"E4",X"02",X"DE",X"C0",X"C0",X"C0",X"C0",X"C0",X"E4",
		X"08",X"DC",X"FC",X"DA",X"02",X"E6",X"E8",X"E8",X"E8",X"E8",X"EA",X"02",X"E7",X"E9",X"E9",X"E9",
		X"E9",X"EB",X"02",X"DE",X"F3",X"E9",X"E9",X"E9",X"E9",X"EB",X"02",X"E6",X"E8",X"E8",X"E8",X"EA",
		X"02",X"DC",X"FC",X"DA",X"02",X"E7",X"E9",X"E9",X"E9",X"F5",X"E4",X"09",X"DE",X"E4",X"07",X"DE",
		X"F3",X"E9",X"E9",X"EB",X"02",X"DC",X"FC",X"DA",X"06",X"DE",X"E4",X"02",X"E6",X"EA",X"02",X"E6",
		X"E8",X"E8",X"E8",X"F4",X"E4",X"02",X"E6",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"05",X"DC",X"FC",
		X"DA",X"02",X"E6",X"E8",X"EA",X"02",X"E7",X"EB",X"02",X"DE",X"E4",X"02",X"E7",X"E9",X"E9",X"E9",
		X"E9",X"EB",X"02",X"E7",X"E9",X"F5",X"E4",X"02",X"E7",X"EB",X"02",X"E6",X"EA",X"02",X"DC",X"FC",
		X"DA",X"02",X"DE",X"C0",X"E4",X"05",X"DE",X"E4",X"0B",X"DE",X"E4",X"05",X"DE",X"E4",X"02",X"DC",
		X"FC",X"DA",X"02",X"DE",X"C0",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"F2",X"E8",X"E8",X"EA",X"02",
		X"E6",X"E8",X"E8",X"E8",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"E4",X"02",X"DC",
		X"FC",X"DA",X"02",X"E7",X"E9",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",X"E9",X"E9",X"E9",X"EB",X"02",
		X"E7",X"E9",X"E9",X"F5",X"E4",X"02",X"E7",X"EB",X"02",X"E7",X"E9",X"E9",X"F5",X"E4",X"02",X"DC",
		X"FC",X"DA",X"12",X"DE",X"E4",X"08",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"E6",X"E8",X"E8",
		X"E8",X"E8",X"EA",X"02",X"E6",X"EA",X"02",X"EC",X"D3",X"D3",X"D3",X"EE",X"02",X"DE",X"E4",X"02",
		X"E6",X"EA",X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"F3",X"E9",
		X"E9",X"E9",X"EB",X"02",X"DE",X"E4",X"02",X"DC",X"04",X"DA",X"02",X"E7",X"EB",X"02",X"DE",X"E4",
		X"02",X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"E4",X"06",X"DE",X"E4",
		X"02",X"DC",X"04",X"DA",X"05",X"DE",X"E4",X"02",X"DE",X"E4",X"05",X"DC",X"FC",X"DA",X"02",X"DE",
		X"E4",X"02",X"E6",X"E8",X"E8",X"E8",X"F4",X"E5",X"02",X"DC",X"04",X"DA",X"02",X"E6",X"E8",X"E8",
		X"F4",X"E4",X"02",X"DE",X"E4",X"02",X"E6",X"E8",X"E8",X"F4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"62",X"01",X"02",X"01",X"01",X"01",X"01",X"0F",X"01",X"01",X"01",X"02",X"01",X"04",X"07",
		X"0F",X"06",X"04",X"07",X"01",X"01",X"01",X"07",X"01",X"01",X"01",X"01",X"01",X"06",X"04",X"01",
		X"01",X"01",X"01",X"03",X"03",X"07",X"05",X"03",X"01",X"01",X"01",X"04",X"04",X"03",X"03",X"07",
		X"05",X"03",X"03",X"04",X"04",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"04",X"04",X"0F",X"03",X"06",X"04",X"04",X"0F",X"03",
		X"06",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0C",X"01",X"01",X"01",X"01",X"01",X"01",
		X"03",X"04",X"07",X"12",X"03",X"04",X"07",X"12",X"03",X"04",X"03",X"01",X"01",X"01",X"01",X"12",
		X"01",X"01",X"01",X"04",X"03",X"16",X"07",X"03",X"16",X"07",X"03",X"01",X"01",X"01",X"01",X"12",
		X"01",X"01",X"01",X"04",X"07",X"12",X"03",X"04",X"07",X"12",X"03",X"04",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"0C",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"04",X"04",X"0F",X"03",X"06",
		X"04",X"04",X"0F",X"03",X"06",X"04",X"04",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"04",X"04",X"03",X"03",X"07",X"05",X"03",
		X"03",X"04",X"01",X"01",X"01",X"01",X"03",X"03",X"07",X"05",X"03",X"01",X"01",X"01",X"04",X"07",
		X"01",X"01",X"01",X"07",X"01",X"01",X"01",X"01",X"01",X"06",X"04",X"07",X"0F",X"06",X"04",X"01",
		X"02",X"01",X"01",X"01",X"01",X"0F",X"01",X"01",X"01",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"A0",
		X"4D",X"A7",X"C8",X"3A",X"AC",X"4D",X"A7",X"C0",X"CD",X"A1",X"1F",X"2A",X"31",X"4D",X"01",X"99",
		X"4D",X"CD",X"27",X"1F",X"3A",X"99",X"4D",X"A7",X"CA",X"62",X"A3",X"2A",X"60",X"4D",X"29",X"22",
		X"60",X"4D",X"2A",X"5E",X"4D",X"ED",X"6A",X"22",X"5E",X"4D",X"D0",X"21",X"60",X"4D",X"34",X"C3",
		X"D0",X"A3",X"3A",X"A7",X"4D",X"A7",X"CA",X"80",X"A3",X"2A",X"5C",X"4D",X"29",X"22",X"5C",X"4D",
		X"2A",X"5A",X"4D",X"ED",X"6A",X"22",X"5A",X"4D",X"D0",X"21",X"5C",X"4D",X"34",X"C3",X"D0",X"A3",
		X"3A",X"B7",X"4D",X"A7",X"CA",X"9E",X"A3",X"2A",X"50",X"4D",X"29",X"22",X"50",X"4D",X"2A",X"4E",
		X"4D",X"ED",X"6A",X"22",X"4E",X"4D",X"D0",X"21",X"50",X"4D",X"34",X"C3",X"D0",X"A3",X"3A",X"B6",
		X"4D",X"A7",X"CA",X"BC",X"A3",X"2A",X"54",X"4D",X"29",X"22",X"54",X"4D",X"2A",X"52",X"4D",X"ED",
		X"6A",X"22",X"52",X"4D",X"D0",X"21",X"54",X"4D",X"34",X"C3",X"D0",X"A3",X"2A",X"58",X"4D",X"29",
		X"22",X"58",X"4D",X"2A",X"56",X"4D",X"ED",X"6A",X"22",X"56",X"4D",X"D0",X"21",X"58",X"4D",X"34",
		X"21",X"14",X"4D",X"7E",X"A7",X"CA",X"E5",X"A3",X"3A",X"00",X"4D",X"E6",X"07",X"FE",X"04",X"CA",
		X"EF",X"A3",X"C3",X"2E",X"A4",X"3A",X"01",X"4D",X"E6",X"07",X"FE",X"04",X"C2",X"2E",X"A4",X"3E",
		X"01",X"CD",X"C8",X"A6",X"38",X"1B",X"3A",X"A7",X"4D",X"A7",X"CA",X"03",X"A4",X"EF",X"0C",X"00",
		X"C3",X"11",X"A4",X"2A",X"0A",X"4D",X"CD",X"1F",X"1F",X"7E",X"FE",X"1A",X"28",X"03",X"EF",X"08",
		X"00",X"CD",X"7D",X"2E",X"DD",X"21",X"1E",X"4D",X"FD",X"21",X"0A",X"4D",X"CD",X"CD",X"1E",X"22",
		X"0A",X"4D",X"2A",X"1E",X"4D",X"22",X"14",X"4D",X"3A",X"2C",X"4D",X"32",X"28",X"4D",X"DD",X"21",
		X"14",X"4D",X"FD",X"21",X"00",X"4D",X"CD",X"CD",X"1E",X"22",X"00",X"4D",X"CD",X"E5",X"1E",X"22",
		X"31",X"4D",X"C9",X"3A",X"A1",X"4D",X"FE",X"01",X"C0",X"3A",X"AD",X"4D",X"A7",X"C0",X"2A",X"33",
		X"4D",X"01",X"9A",X"4D",X"CD",X"27",X"1F",X"3A",X"9A",X"4D",X"A7",X"CA",X"75",X"A4",X"2A",X"6C",
		X"4D",X"29",X"22",X"6C",X"4D",X"2A",X"6A",X"4D",X"ED",X"6A",X"22",X"6A",X"4D",X"D0",X"21",X"6C",
		X"4D",X"34",X"C3",X"A7",X"A4",X"3A",X"A8",X"4D",X"A7",X"CA",X"93",X"A4",X"2A",X"68",X"4D",X"29",
		X"22",X"68",X"4D",X"2A",X"66",X"4D",X"ED",X"6A",X"22",X"66",X"4D",X"D0",X"21",X"68",X"4D",X"34",
		X"C3",X"A7",X"A4",X"2A",X"64",X"4D",X"29",X"22",X"64",X"4D",X"2A",X"62",X"4D",X"ED",X"6A",X"22",
		X"62",X"4D",X"D0",X"21",X"64",X"4D",X"34",X"21",X"16",X"4D",X"7E",X"A7",X"CA",X"BC",X"A4",X"3A",
		X"02",X"4D",X"E6",X"07",X"FE",X"04",X"CA",X"C6",X"A4",X"C3",X"05",X"A5",X"3A",X"03",X"4D",X"E6",
		X"07",X"FE",X"04",X"C2",X"05",X"A5",X"3E",X"02",X"CD",X"C8",X"A6",X"38",X"1B",X"3A",X"A8",X"4D",
		X"A7",X"CA",X"DA",X"A4",X"EF",X"0D",X"00",X"C3",X"E8",X"A4",X"2A",X"0C",X"4D",X"CD",X"1F",X"1F",
		X"7E",X"FE",X"1A",X"28",X"03",X"EF",X"09",X"00",X"CD",X"A4",X"2E",X"DD",X"21",X"20",X"4D",X"FD",
		X"21",X"0C",X"4D",X"CD",X"CD",X"1E",X"22",X"0C",X"4D",X"2A",X"20",X"4D",X"22",X"16",X"4D",X"3A",
		X"2D",X"4D",X"32",X"29",X"4D",X"DD",X"21",X"16",X"4D",X"FD",X"21",X"02",X"4D",X"CD",X"CD",X"1E",
		X"22",X"02",X"4D",X"CD",X"E5",X"1E",X"22",X"33",X"4D",X"C9",X"3A",X"A2",X"4D",X"FE",X"01",X"C0",
		X"3A",X"AE",X"4D",X"A7",X"C0",X"2A",X"35",X"4D",X"01",X"9B",X"4D",X"CD",X"27",X"1F",X"3A",X"9B",
		X"4D",X"A7",X"CA",X"4C",X"A5",X"2A",X"78",X"4D",X"29",X"22",X"78",X"4D",X"2A",X"76",X"4D",X"ED",
		X"6A",X"22",X"76",X"4D",X"D0",X"21",X"78",X"4D",X"34",X"C3",X"7E",X"A5",X"3A",X"A9",X"4D",X"A7",
		X"CA",X"6A",X"A5",X"2A",X"74",X"4D",X"29",X"22",X"74",X"4D",X"2A",X"72",X"4D",X"ED",X"6A",X"22",
		X"72",X"4D",X"D0",X"21",X"74",X"4D",X"34",X"C3",X"7E",X"A5",X"2A",X"70",X"4D",X"29",X"22",X"70",
		X"4D",X"2A",X"6E",X"4D",X"ED",X"6A",X"22",X"6E",X"4D",X"D0",X"21",X"70",X"4D",X"34",X"21",X"18",
		X"4D",X"7E",X"A7",X"CA",X"93",X"A5",X"3A",X"04",X"4D",X"E6",X"07",X"FE",X"04",X"CA",X"9D",X"A5",
		X"C3",X"DC",X"A5",X"3A",X"05",X"4D",X"E6",X"07",X"FE",X"04",X"C2",X"DC",X"A5",X"3E",X"03",X"CD",
		X"C8",X"A6",X"38",X"1B",X"3A",X"A9",X"4D",X"A7",X"CA",X"B1",X"A5",X"EF",X"0E",X"00",X"C3",X"BF",
		X"A5",X"2A",X"0E",X"4D",X"CD",X"1F",X"1F",X"7E",X"FE",X"1A",X"28",X"03",X"EF",X"0A",X"00",X"CD",
		X"CB",X"2E",X"DD",X"21",X"22",X"4D",X"FD",X"21",X"0E",X"4D",X"CD",X"CD",X"1E",X"22",X"0E",X"4D",
		X"2A",X"22",X"4D",X"22",X"18",X"4D",X"3A",X"2E",X"4D",X"32",X"2A",X"4D",X"DD",X"21",X"18",X"4D",
		X"FD",X"21",X"04",X"4D",X"CD",X"CD",X"1E",X"22",X"04",X"4D",X"CD",X"E5",X"1E",X"22",X"35",X"4D",
		X"C9",X"3A",X"A3",X"4D",X"FE",X"01",X"C0",X"3A",X"AF",X"4D",X"A7",X"C0",X"2A",X"37",X"4D",X"01",
		X"9C",X"4D",X"CD",X"27",X"1F",X"3A",X"9C",X"4D",X"A7",X"CA",X"23",X"A6",X"2A",X"84",X"4D",X"29",
		X"22",X"84",X"4D",X"2A",X"82",X"4D",X"ED",X"6A",X"22",X"82",X"4D",X"D0",X"21",X"84",X"4D",X"34",
		X"C3",X"55",X"A6",X"3A",X"AA",X"4D",X"A7",X"CA",X"41",X"A6",X"2A",X"80",X"4D",X"29",X"22",X"80",
		X"4D",X"2A",X"7E",X"4D",X"ED",X"6A",X"22",X"7E",X"4D",X"D0",X"21",X"80",X"4D",X"34",X"C3",X"55",
		X"A6",X"2A",X"7C",X"4D",X"29",X"22",X"7C",X"4D",X"2A",X"7A",X"4D",X"ED",X"6A",X"22",X"7A",X"4D",
		X"D0",X"21",X"7C",X"4D",X"34",X"21",X"1A",X"4D",X"7E",X"A7",X"CA",X"6A",X"A6",X"3A",X"06",X"4D",
		X"E6",X"07",X"FE",X"04",X"CA",X"74",X"A6",X"C3",X"B3",X"A6",X"3A",X"07",X"4D",X"E6",X"07",X"FE",
		X"04",X"C2",X"B3",X"A6",X"3E",X"04",X"CD",X"C8",X"A6",X"38",X"1B",X"3A",X"AA",X"4D",X"A7",X"CA",
		X"88",X"A6",X"EF",X"0F",X"00",X"C3",X"96",X"A6",X"2A",X"10",X"4D",X"CD",X"1F",X"1F",X"7E",X"FE",
		X"1A",X"28",X"03",X"EF",X"0B",X"00",X"CD",X"F2",X"2E",X"DD",X"21",X"24",X"4D",X"FD",X"21",X"10",
		X"4D",X"CD",X"CD",X"1E",X"22",X"10",X"4D",X"2A",X"24",X"4D",X"22",X"1A",X"4D",X"3A",X"2F",X"4D",
		X"32",X"2B",X"4D",X"DD",X"21",X"1A",X"4D",X"FD",X"21",X"06",X"4D",X"CD",X"CD",X"1E",X"22",X"06",
		X"4D",X"CD",X"E5",X"1E",X"22",X"37",X"4D",X"C9",X"87",X"4F",X"06",X"00",X"21",X"09",X"4D",X"09",
		X"7E",X"FE",X"1D",X"C2",X"DB",X"A6",X"36",X"3D",X"C3",X"F4",X"A6",X"FE",X"3E",X"C2",X"E5",X"A6",
		X"36",X"1E",X"C3",X"F4",X"A6",X"06",X"21",X"90",X"DA",X"F4",X"A6",X"7E",X"06",X"3B",X"90",X"D2",
		X"F4",X"A6",X"A7",X"C9",X"37",X"C9",X"41",X"B0",X"41",X"B0",X"37",X"AF",X"C0",X"AC",X"27",X"AC",
		X"86",X"A8",X"84",X"A7",X"86",X"A8",X"C5",X"A9",X"9E",X"AA",X"C5",X"A7",X"14",X"3C",X"3E",X"A8",
		X"C5",X"A9",X"37",X"AF",X"27",X"AC",X"84",X"A7",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",
		X"85",X"A8",X"85",X"A8",X"85",X"A8",X"AA",X"AF",X"AA",X"AF",X"BE",X"AE",X"C0",X"AC",X"8D",X"AC",
		X"26",X"A9",X"A5",X"A7",X"26",X"A9",X"3D",X"AA",X"80",X"AB",X"08",X"A8",X"91",X"3B",X"61",X"A8",
		X"3D",X"AA",X"BE",X"AE",X"8D",X"AC",X"A5",X"A7",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",
		X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"D8",X"AD",X"85",X"A8",X"85",X"A8",X"85",X"A8",
		X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",
		X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",X"85",X"A8",
		X"85",X"A8",X"85",X"A8",X"F1",X"00",X"F2",X"02",X"F3",X"0A",X"F4",X"00",X"41",X"43",X"45",X"86",
		X"8A",X"88",X"8B",X"6A",X"6B",X"71",X"6A",X"88",X"8B",X"6A",X"6B",X"71",X"6A",X"6B",X"71",X"73",
		X"75",X"96",X"95",X"96",X"FF",X"F1",X"02",X"F2",X"03",X"F3",X"0A",X"F4",X"02",X"50",X"70",X"86",
		X"90",X"81",X"90",X"86",X"90",X"68",X"6A",X"6B",X"68",X"6A",X"68",X"66",X"6A",X"68",X"66",X"65",
		X"68",X"86",X"81",X"86",X"FF",X"F1",X"00",X"F2",X"02",X"F3",X"0A",X"F4",X"00",X"69",X"6B",X"69",
		X"86",X"61",X"64",X"65",X"86",X"86",X"64",X"66",X"64",X"61",X"69",X"6B",X"69",X"86",X"61",X"64",
		X"64",X"A1",X"70",X"71",X"74",X"75",X"35",X"76",X"30",X"50",X"35",X"76",X"30",X"50",X"54",X"56",
		X"54",X"51",X"6B",X"69",X"6B",X"69",X"6B",X"91",X"6B",X"69",X"66",X"F2",X"01",X"74",X"76",X"74",
		X"71",X"74",X"71",X"6B",X"69",X"A6",X"A6",X"FF",X"F1",X"03",X"F2",X"03",X"F3",X"0A",X"F4",X"02",
		X"70",X"66",X"70",X"46",X"50",X"86",X"90",X"70",X"66",X"70",X"46",X"50",X"86",X"90",X"70",X"66",
		X"70",X"46",X"50",X"86",X"90",X"70",X"61",X"70",X"41",X"50",X"81",X"90",X"F4",X"00",X"A6",X"A4",
		X"A2",X"A1",X"F4",X"01",X"86",X"89",X"8B",X"81",X"74",X"71",X"6B",X"69",X"A6",X"FF",X"F1",X"00",
		X"F2",X"02",X"F3",X"0A",X"F4",X"00",X"65",X"64",X"65",X"88",X"67",X"88",X"61",X"63",X"64",X"85",
		X"64",X"85",X"6A",X"69",X"6A",X"8C",X"75",X"93",X"90",X"91",X"90",X"91",X"70",X"8A",X"68",X"71",
		X"FF",X"F1",X"02",X"F2",X"03",X"F3",X"0A",X"F4",X"02",X"65",X"90",X"68",X"70",X"68",X"67",X"66",
		X"65",X"90",X"61",X"70",X"61",X"65",X"68",X"66",X"90",X"63",X"90",X"86",X"90",X"85",X"90",X"85",
		X"70",X"86",X"68",X"65",X"FF",X"FF",X"F1",X"00",X"F2",X"01",X"F3",X"0A",X"F4",X"00",X"77",X"76",
		X"57",X"50",X"97",X"F2",X"02",X"74",X"92",X"8C",X"F2",X"01",X"90",X"90",X"90",X"74",X"73",X"74",
		X"75",X"77",X"75",X"74",X"72",X"74",X"73",X"74",X"8C",X"67",X"6C",X"72",X"74",X"73",X"74",X"75",
		X"77",X"7C",X"7B",X"79",X"77",X"75",X"72",X"6B",X"8B",X"90",X"77",X"75",X"72",X"8B",X"6C",X"6E",
		X"6F",X"74",X"75",X"76",X"97",X"70",X"7C",X"70",X"7B",X"77",X"74",X"6C",X"6B",X"73",X"76",X"77",
		X"94",X"74",X"76",X"77",X"70",X"74",X"70",X"7B",X"70",X"79",X"70",X"77",X"70",X"76",X"70",X"F2",
		X"02",X"74",X"73",X"74",X"6B",X"6B",X"6A",X"6B",X"67",X"F2",X"01",X"77",X"76",X"77",X"74",X"74",
		X"70",X"74",X"70",X"73",X"74",X"76",X"77",X"79",X"7C",X"7B",X"59",X"50",X"79",X"77",X"76",X"97",
		X"70",X"74",X"70",X"F2",X"02",X"74",X"F2",X"01",X"7C",X"79",X"76",X"56",X"50",X"76",X"79",X"5C",
		X"50",X"7C",X"7B",X"7A",X"9B",X"70",X"74",X"70",X"73",X"74",X"76",X"77",X"79",X"7C",X"7B",X"73",
		X"94",X"91",X"F2",X"02",X"74",X"FF",X"F1",X"03",X"F2",X"03",X"F3",X"06",X"F4",X"03",X"87",X"90",
		X"87",X"90",X"6C",X"70",X"67",X"70",X"69",X"70",X"6B",X"70",X"6C",X"70",X"74",X"70",X"67",X"70",
		X"6B",X"70",X"6C",X"70",X"74",X"70",X"67",X"70",X"74",X"70",X"6C",X"70",X"77",X"70",X"74",X"70",
		X"73",X"70",X"72",X"70",X"77",X"70",X"67",X"70",X"75",X"70",X"6B",X"70",X"75",X"70",X"67",X"70",
		X"6B",X"70",X"6C",X"70",X"77",X"70",X"74",X"70",X"77",X"70",X"6B",X"70",X"7B",X"70",X"6B",X"70",
		X"7B",X"70",X"F4",X"00",X"94",X"74",X"76",X"77",X"F4",X"01",X"70",X"74",X"70",X"6B",X"70",X"6C",
		X"70",X"6D",X"70",X"6F",X"70",X"74",X"70",X"77",X"70",X"6B",X"70",X"74",X"70",X"F3",X"0A",X"67",
		X"70",X"6B",X"70",X"64",X"70",X"67",X"70",X"66",X"70",X"6F",X"70",X"6B",X"70",X"6F",X"70",X"64",
		X"70",X"6B",X"70",X"67",X"70",X"74",X"70",X"69",X"70",X"76",X"70",X"6B",X"70",X"6F",X"70",X"64",
		X"70",X"6B",X"70",X"67",X"70",X"77",X"70",X"6B",X"70",X"7B",X"70",X"6B",X"70",X"7B",X"70",X"74",
		X"70",X"6B",X"70",X"64",X"FF",X"F1",X"00",X"F2",X"02",X"F3",X"08",X"F4",X"01",X"B0",X"B0",X"90",
		X"74",X"74",X"73",X"74",X"F4",X"00",X"97",X"77",X"94",X"74",X"F4",X"01",X"87",X"67",X"93",X"72",
		X"8C",X"90",X"90",X"87",X"74",X"74",X"73",X"74",X"F4",X"00",X"8C",X"6C",X"97",X"77",X"F4",X"01",
		X"95",X"74",X"92",X"74",X"F4",X"00",X"95",X"75",X"90",X"70",X"F4",X"01",X"79",X"78",X"79",X"75",
		X"74",X"75",X"F4",X"00",X"92",X"72",X"97",X"77",X"F4",X"01",X"94",X"73",X"94",X"75",X"97",X"75",
		X"94",X"72",X"87",X"74",X"74",X"73",X"74",X"F4",X"00",X"97",X"77",X"94",X"74",X"F4",X"01",X"96",
		X"76",X"76",X"74",X"76",X"F4",X"00",X"99",X"79",X"90",X"79",X"F4",X"01",X"77",X"76",X"74",X"9B",
		X"74",X"73",X"71",X"6B",X"96",X"77",X"F4",X"00",X"94",X"94",X"94",X"94",X"FF",X"F1",X"03",X"F2",
		X"03",X"F3",X"08",X"F4",X"00",X"B0",X"B0",X"8C",X"6C",X"94",X"74",X"97",X"F4",X"01",X"6C",X"6C",
		X"6B",X"6C",X"87",X"F4",X"00",X"67",X"89",X"6B",X"8C",X"67",X"89",X"6B",X"8C",X"74",X"87",X"74",
		X"8C",X"74",X"87",X"74",X"92",X"75",X"87",X"75",X"8B",X"75",X"87",X"75",X"8B",X"75",X"87",X"75",
		X"8B",X"75",X"87",X"72",X"8C",X"74",X"87",X"74",X"8B",X"67",X"89",X"6B",X"8C",X"74",X"87",X"74",
		X"8C",X"74",X"87",X"74",X"8B",X"73",X"86",X"73",X"F4",X"01",X"8B",X"6B",X"F4",X"00",X"91",X"73",
		X"94",X"94",X"70",X"74",X"8B",X"8B",X"60",X"6B",X"94",X"6B",X"87",X"6B",X"84",X"FF",X"F1",X"00",
		X"F2",X"02",X"F3",X"0A",X"F4",X"00",X"59",X"58",X"59",X"50",X"54",X"53",X"54",X"50",X"4C",X"4B",
		X"4C",X"50",X"49",X"48",X"49",X"50",X"44",X"43",X"24",X"30",X"64",X"4C",X"6B",X"89",X"69",X"70",
		X"59",X"58",X"59",X"50",X"59",X"58",X"59",X"50",X"59",X"58",X"59",X"74",X"50",X"74",X"55",X"54",
		X"55",X"50",X"59",X"58",X"59",X"50",X"94",X"74",X"6C",X"52",X"51",X"52",X"50",X"4B",X"4A",X"4B",
		X"50",X"55",X"54",X"55",X"68",X"48",X"72",X"4C",X"4B",X"4C",X"50",X"46",X"44",X"46",X"50",X"88",
		X"68",X"64",X"59",X"58",X"59",X"50",X"59",X"58",X"59",X"50",X"59",X"58",X"59",X"74",X"54",X"77",
		X"55",X"54",X"55",X"50",X"4C",X"4B",X"4C",X"50",X"95",X"75",X"76",X"57",X"56",X"57",X"50",X"47",
		X"46",X"47",X"50",X"57",X"56",X"57",X"50",X"5C",X"5B",X"5C",X"50",X"47",X"46",X"27",X"30",X"67",
		X"54",X"72",X"8C",X"6C",X"67",X"54",X"53",X"74",X"4C",X"4B",X"6C",X"54",X"53",X"54",X"77",X"59",
		X"77",X"55",X"54",X"75",X"4B",X"49",X"6B",X"95",X"75",X"70",X"47",X"46",X"67",X"4B",X"4A",X"6B",
		X"59",X"58",X"59",X"4B",X"6B",X"57",X"50",X"57",X"59",X"57",X"50",X"57",X"59",X"57",X"50",X"77",
		X"75",X"74",X"72",X"54",X"53",X"74",X"4C",X"4B",X"6C",X"57",X"56",X"57",X"54",X"74",X"77",X"59",
		X"58",X"59",X"50",X"59",X"58",X"59",X"3C",X"30",X"9C",X"7C",X"79",X"57",X"59",X"77",X"54",X"55",
		X"74",X"4C",X"4E",X"4C",X"47",X"67",X"77",X"47",X"46",X"27",X"30",X"67",X"54",X"72",X"AC",X"FF",
		X"F1",X"03",X"F2",X"03",X"F3",X"08",X"F4",X"02",X"79",X"70",X"74",X"70",X"6C",X"70",X"69",X"70",
		X"64",X"70",X"64",X"70",X"69",X"6C",X"64",X"6C",X"69",X"74",X"64",X"74",X"69",X"74",X"64",X"74",
		X"6B",X"72",X"64",X"72",X"69",X"6C",X"64",X"74",X"6B",X"74",X"64",X"74",X"68",X"72",X"64",X"6B",
		X"69",X"74",X"62",X"6C",X"64",X"74",X"64",X"74",X"69",X"74",X"64",X"74",X"69",X"74",X"64",X"74",
		X"65",X"6C",X"F2",X"02",X"60",X"F2",X"03",X"6C",X"65",X"6C",X"F2",X"02",X"60",X"F2",X"03",X"6C",
		X"6C",X"74",X"67",X"6C",X"64",X"67",X"F2",X"02",X"60",X"F2",X"03",X"6C",X"67",X"77",X"67",X"77",
		X"F2",X"01",X"7C",X"F2",X"03",X"6C",X"6C",X"5C",X"50",X"F2",X"04",X"6C",X"74",X"67",X"74",X"6C",
		X"74",X"67",X"74",X"6B",X"75",X"67",X"75",X"6B",X"75",X"67",X"75",X"6B",X"75",X"67",X"75",X"6B",
		X"75",X"67",X"6B",X"6C",X"74",X"67",X"74",X"6B",X"67",X"69",X"6B",X"6C",X"74",X"67",X"74",X"6C",
		X"74",X"67",X"74",X"65",X"6C",X"F2",X"02",X"60",X"F2",X"04",X"6C",X"65",X"6C",X"69",X"66",X"67",
		X"74",X"6C",X"74",X"67",X"74",X"6C",X"FF",X"F1",X"00",X"F2",X"02",X"F3",X"0A",X"F4",X"06",X"B5",
		X"96",X"98",X"98",X"96",X"95",X"93",X"91",X"91",X"93",X"95",X"95",X"F5",X"73",X"B3",X"B5",X"96",
		X"98",X"98",X"96",X"95",X"93",X"91",X"91",X"93",X"95",X"93",X"F5",X"71",X"B1",X"B3",X"95",X"91",
		X"93",X"75",X"76",X"95",X"91",X"93",X"75",X"76",X"95",X"93",X"91",X"93",X"88",X"B5",X"90",X"96",
		X"98",X"98",X"96",X"95",X"93",X"91",X"91",X"93",X"95",X"93",X"F5",X"71",X"B1",X"B3",X"95",X"91",
		X"93",X"75",X"76",X"95",X"91",X"93",X"75",X"76",X"95",X"93",X"91",X"93",X"88",X"B5",X"90",X"96",
		X"98",X"98",X"96",X"95",X"93",X"91",X"91",X"93",X"95",X"93",X"71",X"B1",X"FF",X"F1",X"02",X"F2",
		X"03",X"F3",X"08",X"F4",X"06",X"D1",X"C8",X"D1",X"C8",X"D1",X"C8",X"D1",X"A8",X"B1",X"B8",X"B1",
		X"B8",X"B1",X"F2",X"04",X"A3",X"A5",X"F2",X"03",X"BA",X"93",X"98",X"D1",X"C8",X"D1",X"A8",X"B1",
		X"B8",X"B1",X"B8",X"B1",X"B3",X"B5",X"AA",X"93",X"98",X"D1",X"C8",X"D1",X"A8",X"B1",X"FF",X"FF",
		X"F1",X"03",X"F2",X"04",X"F3",X"0A",X"F4",X"06",X"49",X"8A",X"70",X"F5",X"4C",X"91",X"70",X"F5",
		X"49",X"6A",X"F5",X"4C",X"71",X"F5",X"56",X"75",X"F5",X"4A",X"71",X"F5",X"55",X"B4",X"75",X"73",
		X"71",X"6A",X"68",X"AA",X"F5",X"70",X"F5",X"49",X"8A",X"70",X"F5",X"4C",X"91",X"70",X"F5",X"48",
		X"6A",X"F5",X"4C",X"61",X"F5",X"56",X"75",X"F5",X"51",X"75",X"F5",X"5A",X"D9",X"B9",X"F5",X"70",
		X"F5",X"49",X"8A",X"70",X"F5",X"4C",X"91",X"70",X"F5",X"49",X"6A",X"F5",X"4C",X"71",X"F5",X"56",
		X"75",X"F5",X"4A",X"71",X"F5",X"55",X"B4",X"75",X"73",X"71",X"6A",X"68",X"6A",X"CA",X"90",X"7A",
		X"F5",X"58",X"75",X"F5",X"53",X"71",X"F5",X"4A",X"54",X"73",X"F5",X"55",X"73",X"F5",X"55",X"73",
		X"F5",X"55",X"73",X"F5",X"71",X"6A",X"68",X"6A",X"6A",X"AA",X"AA",X"F5",X"90",X"71",X"6A",X"68",
		X"6A",X"6A",X"AA",X"AA",X"F5",X"90",X"71",X"6A",X"68",X"6A",X"6A",X"AA",X"AA",X"F5",X"70",X"F5",
		X"89",X"8A",X"70",X"F5",X"4C",X"91",X"70",X"F5",X"49",X"6A",X"F5",X"4C",X"71",X"F5",X"56",X"75",
		X"F5",X"4A",X"71",X"F5",X"55",X"B4",X"75",X"73",X"71",X"6A",X"68",X"AA",X"F5",X"70",X"F5",X"49",
		X"8A",X"70",X"F5",X"4C",X"91",X"70",X"F5",X"48",X"6A",X"F5",X"4C",X"61",X"F5",X"56",X"75",X"F5",
		X"51",X"75",X"F5",X"5A",X"D9",X"B9",X"F5",X"70",X"F5",X"49",X"8A",X"70",X"F5",X"4C",X"91",X"70",
		X"F5",X"49",X"6A",X"F5",X"4C",X"71",X"F5",X"56",X"75",X"F5",X"4A",X"71",X"F5",X"55",X"B4",X"75",
		X"73",X"71",X"6A",X"68",X"6A",X"CA",X"90",X"7A",X"F5",X"58",X"75",X"F5",X"53",X"71",X"F5",X"4A",
		X"54",X"73",X"F5",X"55",X"73",X"F5",X"55",X"73",X"F5",X"55",X"73",X"F5",X"71",X"6A",X"68",X"6A",
		X"6A",X"AA",X"AA",X"F5",X"90",X"71",X"6A",X"68",X"6A",X"6A",X"AA",X"AA",X"F5",X"90",X"71",X"6A",
		X"68",X"6A",X"6A",X"AA",X"AA",X"F5",X"90",X"FF",X"F1",X"00",X"F2",X"01",X"F3",X"08",X"F4",X"00",
		X"B5",X"B5",X"B3",X"B3",X"71",X"6C",X"71",X"73",X"71",X"6A",X"65",X"66",X"68",X"6A",X"68",X"3E",
		X"43",X"3E",X"11",X"3E",X"2F",X"6F",X"3E",X"42",X"3E",X"42",X"3E",X"42",X"67",X"7E",X"FE",X"4D",
		X"20",X"ED",X"19",X"6F",X"3E",X"42",X"67",X"3E",X"42",X"FE",X"4D",X"FE",X"4D",X"FE",X"4D",X"7E",
		X"E1",X"E9",X"9D",X"9D",X"98",X"98",X"95",X"95",X"93",X"71",X"73",X"95",X"98",X"78",X"75",X"71",
		X"FF",X"F1",X"00",X"F2",X"01",X"F3",X"08",X"F4",X"00",X"B5",X"B5",X"B3",X"B3",X"71",X"6C",X"71",
		X"73",X"71",X"6A",X"65",X"66",X"68",X"6A",X"68",X"01",X"00",X"40",X"DD",X"21",X"00",X"00",X"21",
		X"00",X"00",X"16",X"00",X"7E",X"5F",X"DD",X"19",X"32",X"C0",X"50",X"23",X"0B",X"79",X"B0",X"20",
		X"F1",X"11",X"00",X"40",X"19",X"01",X"00",X"40",X"16",X"00",X"7E",X"5F",X"DD",X"19",X"32",X"C0",
		X"50",X"23",X"0B",X"79",X"B0",X"20",X"F1",X"DD",X"E5",X"E1",X"7D",X"AF",X"C9",X"08",X"3A",X"00",
		X"50",X"CB",X"67",X"C2",X"54",X"BC",X"3A",X"00",X"50",X"E6",X"E0",X"FE",X"E0",X"21",X"21",X"C3",
		X"E5",X"C8",X"CD",X"41",X"25",X"08",X"F5",X"DD",X"21",X"50",X"40",X"CD",X"BF",X"24",X"F1",X"47",
		X"AF",X"90",X"DD",X"21",X"55",X"40",X"CD",X"BF",X"24",X"06",X"80",X"CD",X"79",X"32",X"C9",X"E9",
		X"E9",X"E9",X"E9",X"E9",X"C8",X"C8",X"9D",X"9D",X"98",X"98",X"95",X"95",X"93",X"71",X"73",X"95",
		X"98",X"78",X"75",X"71",X"FF",X"F1",X"00",X"F2",X"00",X"F3",X"00",X"F4",X"00",X"FF",X"F1",X"03",
		X"F2",X"03",X"F3",X"06",X"F4",X"03",X"B5",X"B5",X"B3",X"B3",X"91",X"9F",X"88",X"9F",X"91",X"9F",
		X"88",X"9F",X"91",X"9F",X"88",X"9F",X"88",X"9F",X"88",X"9F",X"91",X"9F",X"88",X"9F",X"91",X"9F",
		X"88",X"9F",X"91",X"9F",X"88",X"9F",X"91",X"9F",X"7F",X"7F",X"7D",X"7F",X"7D",X"7C",X"7A",X"78",
		X"7A",X"78",X"76",X"75",X"78",X"76",X"75",X"73",X"51",X"52",X"53",X"54",X"55",X"56",X"78",X"76",
		X"78",X"7A",X"7D",X"7A",X"7C",X"7D",X"7F",X"F2",X"04",X"61",X"63",X"65",X"66",X"F2",X"03",X"46",
		X"4A",X"51",X"53",X"56",X"58",X"5A",X"5D",X"91",X"9F",X"93",X"9F",X"95",X"9F",X"88",X"9F",X"91",
		X"9F",X"88",X"9F",X"91",X"9F",X"98",X"75",X"73",X"F0",X"26",X"A9",X"FF",X"C3",X"EF",X"BF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"00",X"F2",X"01",X"F3",X"08",X"F4",X"00",X"B5",
		X"B5",X"B3",X"B3",X"71",X"6C",X"71",X"73",X"71",X"6A",X"65",X"66",X"68",X"6A",X"68",X"65",X"88",
		X"71",X"73",X"95",X"95",X"75",X"73",X"71",X"73",X"75",X"73",X"73",X"72",X"93",X"75",X"73",X"71",
		X"6C",X"71",X"73",X"71",X"6A",X"65",X"66",X"68",X"6A",X"68",X"65",X"88",X"71",X"73",X"95",X"98",
		X"78",X"76",X"71",X"73",X"75",X"71",X"93",X"B1",X"75",X"98",X"75",X"98",X"98",X"75",X"98",X"75",
		X"58",X"46",X"48",X"4C",X"51",X"55",X"58",X"55",X"76",X"9A",X"76",X"9A",X"9A",X"76",X"9A",X"76",
		X"9A",X"6A",X"6C",X"9D",X"9D",X"98",X"98",X"95",X"95",X"93",X"71",X"73",X"95",X"98",X"78",X"75",
		X"71",X"73",X"75",X"71",X"93",X"B1",X"F0",X"86",X"A8",X"FF",X"F1",X"03",X"F2",X"03",X"F3",X"08",
		X"F4",X"06",X"8A",X"9A",X"8A",X"9A",X"8A",X"9A",X"8A",X"9A",X"83",X"93",X"83",X"93",X"88",X"98",
		X"88",X"98",X"81",X"91",X"81",X"91",X"81",X"91",X"81",X"91",X"8A",X"9A",X"8A",X"9A",X"8A",X"9A",
		X"8A",X"9A",X"83",X"93",X"83",X"93",X"88",X"98",X"88",X"98",X"81",X"91",X"81",X"91",X"81",X"91",
		X"81",X"91",X"83",X"93",X"83",X"93",X"83",X"93",X"83",X"93",X"83",X"93",X"83",X"93",X"83",X"93",
		X"A6",X"A8",X"A8",X"88",X"98",X"88",X"98",X"D5",X"D0",X"8A",X"9A",X"8A",X"9A",X"8A",X"9A",X"8A",
		X"9A",X"83",X"93",X"83",X"93",X"88",X"98",X"88",X"98",X"81",X"91",X"81",X"91",X"81",X"91",X"81",
		X"91",X"8A",X"9A",X"8A",X"9A",X"8A",X"9A",X"8A",X"9A",X"83",X"93",X"83",X"93",X"88",X"98",X"88",
		X"98",X"81",X"91",X"81",X"91",X"81",X"91",X"81",X"91",X"83",X"93",X"83",X"93",X"83",X"93",X"83",
		X"93",X"83",X"93",X"83",X"93",X"83",X"93",X"A6",X"A8",X"A8",X"88",X"98",X"88",X"98",X"D5",X"D0",
		X"FF",X"F1",X"00",X"F2",X"01",X"F3",X"04",X"F4",X"06",X"D5",X"93",X"91",X"8C",X"8A",X"8A",X"91",
		X"8C",X"8A",X"88",X"8A",X"88",X"85",X"C8",X"D0",X"D5",X"93",X"91",X"8C",X"8A",X"8A",X"91",X"8C",
		X"8A",X"88",X"8A",X"88",X"85",X"C8",X"D0",X"93",X"93",X"93",X"91",X"A6",X"86",X"8A",X"95",X"95",
		X"95",X"93",X"A6",X"8A",X"91",X"91",X"F5",X"6A",X"88",X"88",X"88",X"8A",X"88",X"CA",X"D0",X"D5",
		X"93",X"91",X"8C",X"8A",X"8A",X"91",X"8C",X"8A",X"88",X"8A",X"88",X"85",X"C8",X"D0",X"D5",X"93",
		X"91",X"8C",X"8A",X"8A",X"91",X"8C",X"8A",X"88",X"8A",X"88",X"85",X"A8",X"B0",X"93",X"93",X"93",
		X"91",X"A6",X"86",X"8A",X"95",X"95",X"95",X"93",X"A6",X"8A",X"91",X"91",X"F5",X"6A",X"88",X"88",
		X"88",X"8A",X"88",X"CA",X"D0",X"FF",X"2A",X"0A",X"4C",X"22",X"C2",X"4F",X"2A",X"0C",X"4C",X"22",
		X"D3",X"4F",X"2A",X"08",X"4D",X"22",X"C4",X"4F",X"2A",X"D2",X"4D",X"22",X"D0",X"4F",X"2A",X"1A",
		X"4C",X"22",X"D5",X"4F",X"2A",X"1C",X"4C",X"22",X"D7",X"4F",X"C9",X"2A",X"C2",X"4F",X"3E",X"09",
		X"67",X"22",X"0A",X"4C",X"2A",X"D3",X"4F",X"3E",X"05",X"67",X"22",X"0C",X"4C",X"2A",X"C4",X"4F",
		X"22",X"08",X"4D",X"2A",X"D0",X"4F",X"22",X"D2",X"4D",X"2A",X"D5",X"4F",X"22",X"1A",X"4C",X"2A",
		X"D7",X"4F",X"22",X"1C",X"4C",X"C9",X"2A",X"D3",X"4F",X"22",X"0A",X"4C",X"2A",X"D0",X"4F",X"22",
		X"08",X"4D",X"2A",X"D7",X"4F",X"22",X"1A",X"4C",X"C9",X"2A",X"0A",X"4C",X"22",X"D3",X"4F",X"2A",
		X"08",X"4D",X"22",X"D0",X"4F",X"2A",X"1A",X"4C",X"22",X"D7",X"4F",X"C9",X"C9",X"F5",X"2A",X"12",
		X"4D",X"E5",X"2A",X"C6",X"4F",X"22",X"12",X"4D",X"E1",X"22",X"C6",X"4F",X"2A",X"39",X"4D",X"E5",
		X"2A",X"C8",X"4F",X"22",X"39",X"4D",X"E1",X"22",X"C8",X"4F",X"2A",X"1C",X"4D",X"E5",X"2A",X"CA",
		X"4F",X"22",X"1C",X"4D",X"E1",X"22",X"CA",X"4F",X"2A",X"26",X"4D",X"E5",X"2A",X"CC",X"4F",X"22",
		X"26",X"4D",X"E1",X"22",X"CC",X"4F",X"3A",X"30",X"4D",X"F5",X"3A",X"CE",X"4F",X"32",X"30",X"4D",
		X"F1",X"32",X"CE",X"4F",X"3A",X"3C",X"4D",X"F5",X"3A",X"CF",X"4F",X"32",X"3C",X"4D",X"F1",X"32",
		X"CF",X"4F",X"F1",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"98",X"B1",X"FD",
		X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"C9",X"AF",X"32",X"04",X"50",X"32",X"05",X"50",X"3E",
		X"01",X"32",X"00",X"4F",X"3A",X"E0",X"4D",X"FE",X"0F",X"C4",X"04",X"97",X"3A",X"E0",X"4D",X"E7",
		X"C8",X"B1",X"FB",X"B1",X"05",X"B2",X"0F",X"B2",X"19",X"B2",X"23",X"B2",X"2D",X"B2",X"37",X"B2",
		X"41",X"B2",X"4B",X"B2",X"55",X"B2",X"DC",X"B2",X"EF",X"00",X"01",X"EF",X"01",X"00",X"EF",X"04",
		X"00",X"EF",X"1E",X"00",X"21",X"84",X"36",X"11",X"E8",X"4D",X"01",X"10",X"00",X"77",X"ED",X"B0",
		X"EF",X"1C",X"00",X"0E",X"0C",X"06",X"1C",X"CD",X"42",X"00",X"0E",X"0F",X"06",X"20",X"CD",X"42",
		X"00",X"3E",X"27",X"32",X"04",X"4E",X"21",X"E0",X"4D",X"34",X"C9",X"EF",X"20",X"26",X"DD",X"21",
		X"EA",X"4D",X"C3",X"5F",X"B2",X"EF",X"20",X"27",X"DD",X"21",X"EB",X"4D",X"C3",X"5F",X"B2",X"EF",
		X"20",X"28",X"DD",X"21",X"EC",X"4D",X"C3",X"5F",X"B2",X"EF",X"20",X"29",X"DD",X"21",X"ED",X"4D",
		X"C3",X"5F",X"B2",X"EF",X"20",X"2A",X"DD",X"21",X"EE",X"4D",X"C3",X"5F",X"B2",X"EF",X"20",X"2B",
		X"DD",X"21",X"EF",X"4D",X"C3",X"5F",X"B2",X"EF",X"20",X"2C",X"DD",X"21",X"F0",X"4D",X"C3",X"5F",
		X"B2",X"EF",X"20",X"2D",X"DD",X"21",X"F1",X"4D",X"C3",X"5F",X"B2",X"EF",X"20",X"2E",X"DD",X"21",
		X"F2",X"4D",X"C3",X"5F",X"B2",X"EF",X"20",X"2F",X"DD",X"21",X"F3",X"4D",X"C3",X"5F",X"B2",X"3A",
		X"E1",X"4D",X"57",X"3A",X"00",X"50",X"4F",X"32",X"E1",X"4D",X"B2",X"A9",X"32",X"E2",X"4D",X"CB",
		X"57",X"20",X"19",X"CB",X"4F",X"20",X"3D",X"CB",X"5F",X"3E",X"27",X"32",X"04",X"4E",X"C8",X"EF",
		X"1C",X"00",X"21",X"E0",X"4D",X"34",X"3E",X"27",X"32",X"04",X"4E",X"C9",X"DD",X"7E",X"00",X"3C",
		X"FE",X"5A",X"30",X"0F",X"DD",X"77",X"00",X"32",X"02",X"4F",X"EF",X"1C",X"00",X"3E",X"27",X"32",
		X"04",X"4E",X"C9",X"3E",X"5A",X"32",X"02",X"4F",X"DD",X"77",X"00",X"EF",X"1C",X"00",X"3E",X"27",
		X"32",X"04",X"4E",X"C9",X"DD",X"7E",X"00",X"3D",X"FE",X"40",X"38",X"0F",X"32",X"02",X"4F",X"DD",
		X"77",X"00",X"EF",X"1C",X"00",X"3E",X"27",X"32",X"04",X"4E",X"C9",X"3E",X"40",X"32",X"02",X"4F",
		X"DD",X"77",X"00",X"EF",X"1C",X"00",X"3E",X"27",X"32",X"04",X"4E",X"C9",X"21",X"D4",X"83",X"22",
		X"E8",X"4D",X"EF",X"1C",X"00",X"AF",X"32",X"E0",X"4D",X"3A",X"FF",X"4D",X"32",X"04",X"4E",X"AF",
		X"32",X"00",X"4F",X"32",X"00",X"4F",X"32",X"FE",X"4D",X"C9",X"3E",X"40",X"67",X"AF",X"6F",X"3E",
		X"C9",X"77",X"3A",X"70",X"4C",X"FE",X"03",X"C0",X"3A",X"0E",X"4E",X"FE",X"80",X"D8",X"DD",X"2A",
		X"00",X"4C",X"3E",X"1C",X"DD",X"BE",X"02",X"CA",X"90",X"B3",X"DD",X"BE",X"04",X"CA",X"90",X"B3",
		X"DD",X"BE",X"06",X"CA",X"90",X"B3",X"DD",X"BE",X"08",X"CA",X"90",X"B3",X"3A",X"0E",X"4E",X"E6",
		X"01",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"47",X"3A",X"05",X"4E",X"3C",X"80",X"32",X"05",X"4E",
		X"E6",X"7F",X"FE",X"40",X"38",X"02",X"18",X"48",X"DD",X"2A",X"00",X"4C",X"3E",X"1C",X"DD",X"BE",
		X"02",X"C8",X"DD",X"BE",X"04",X"C8",X"DD",X"BE",X"06",X"C8",X"DD",X"BE",X"08",X"C8",X"2A",X"FB",
		X"4D",X"7C",X"B5",X"C0",X"3A",X"FD",X"4D",X"FE",X"05",X"C8",X"21",X"35",X"95",X"CD",X"A1",X"94",
		X"69",X"60",X"3A",X"08",X"4D",X"47",X"3A",X"FD",X"4D",X"80",X"E6",X"03",X"CB",X"27",X"5F",X"16",
		X"00",X"19",X"5E",X"23",X"56",X"EB",X"22",X"FB",X"4D",X"CD",X"1E",X"B4",X"CD",X"A6",X"3F",X"C9",
		X"2A",X"FB",X"4D",X"7C",X"B5",X"C8",X"CD",X"39",X"B4",X"21",X"00",X"00",X"22",X"FB",X"4D",X"C9",
		X"E5",X"21",X"76",X"3A",X"3A",X"13",X"4E",X"E6",X"07",X"CB",X"27",X"5F",X"16",X"00",X"19",X"EB",
		X"E1",X"CD",X"ED",X"B3",X"C9",X"21",X"40",X"86",X"3A",X"13",X"4E",X"78",X"3A",X"08",X"4D",X"81",
		X"83",X"82",X"80",X"ED",X"44",X"E6",X"07",X"CB",X"27",X"5F",X"16",X"00",X"19",X"C9",X"DD",X"E5",
		X"DD",X"21",X"02",X"4C",X"06",X"04",X"CD",X"B5",X"B3",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",
		X"77",X"01",X"DD",X"23",X"DD",X"23",X"10",X"EE",X"DD",X"E1",X"C3",X"58",X"1E",X"1A",X"CD",X"0A",
		X"B4",X"3E",X"04",X"84",X"67",X"13",X"1A",X"CD",X"FB",X"B3",X"C9",X"E5",X"D5",X"77",X"23",X"77",
		X"11",X"1F",X"00",X"19",X"77",X"23",X"77",X"D1",X"E1",X"C9",X"E5",X"D5",X"11",X"1F",X"00",X"77",
		X"3C",X"3C",X"23",X"77",X"3D",X"19",X"77",X"3C",X"3C",X"23",X"77",X"D1",X"E1",X"C9",X"E5",X"D5",
		X"11",X"1F",X"00",X"7E",X"32",X"E3",X"4D",X"23",X"7E",X"32",X"E4",X"4D",X"19",X"7E",X"32",X"E5",
		X"4D",X"23",X"7E",X"32",X"E6",X"4D",X"D1",X"E1",X"C9",X"E5",X"D5",X"11",X"1F",X"00",X"3A",X"E3",
		X"4D",X"77",X"23",X"3A",X"E4",X"4D",X"77",X"19",X"3A",X"E5",X"4D",X"77",X"23",X"3A",X"E6",X"4D",
		X"77",X"D1",X"E1",X"E5",X"D5",X"3E",X"04",X"84",X"67",X"3A",X"7E",X"44",X"77",X"23",X"77",X"11",
		X"1F",X"00",X"19",X"77",X"23",X"77",X"D1",X"E1",X"C9",X"3A",X"13",X"4E",X"3A",X"02",X"4D",X"80",
		X"99",X"82",X"0F",X"0F",X"0F",X"85",X"6F",X"3A",X"00",X"4D",X"85",X"6F",X"3A",X"04",X"4D",X"85",
		X"6F",X"3A",X"06",X"4D",X"85",X"E6",X"0F",X"E7",X"EF",X"B5",X"EF",X"B5",X"FD",X"B5",X"0B",X"B6",
		X"19",X"B6",X"27",X"B6",X"35",X"B6",X"43",X"B6",X"27",X"B6",X"27",X"B6",X"43",X"B6",X"27",X"B6",
		X"35",X"B6",X"43",X"B6",X"43",X"B6",X"51",X"B6",X"51",X"B6",X"51",X"B6",X"1D",X"03",X"5C",X"40",
		X"4F",X"4A",X"45",X"44",X"41",X"40",X"31",X"39",X"39",X"30",X"2F",X"81",X"2F",X"80",X"45",X"03",
		X"40",X"26",X"40",X"40",X"44",X"4F",X"42",X"4C",X"45",X"40",X"40",X"43",X"4F",X"4D",X"41",X"4E",
		X"44",X"4F",X"40",X"40",X"27",X"40",X"2F",X"80",X"2F",X"80",X"45",X"03",X"40",X"26",X"40",X"40",
		X"44",X"4F",X"42",X"4C",X"45",X"40",X"40",X"43",X"4F",X"4D",X"41",X"4E",X"44",X"4F",X"40",X"40",
		X"27",X"40",X"2F",X"81",X"2F",X"80",X"92",X"02",X"40",X"40",X"54",X"55",X"52",X"42",X"4F",X"5B",
		X"40",X"40",X"2F",X"81",X"2F",X"80",X"92",X"02",X"45",X"58",X"54",X"52",X"41",X"40",X"43",X"4F",
		X"49",X"4E",X"2F",X"89",X"2F",X"80",X"9B",X"02",X"4D",X"49",X"4B",X"59",X"40",X"40",X"53",X"52",
		X"4C",X"2F",X"89",X"2F",X"80",X"9B",X"02",X"4D",X"49",X"4B",X"59",X"40",X"40",X"53",X"52",X"4C",
		X"2F",X"81",X"2F",X"80",X"8B",X"02",X"40",X"40",X"4C",X"41",X"4D",X"42",X"41",X"44",X"41",X"2F",
		X"85",X"2F",X"80",X"8E",X"02",X"42",X"55",X"55",X"55",X"55",X"5B",X"40",X"2F",X"8F",X"2F",X"80",
		X"10",X"02",X"4A",X"49",X"40",X"4A",X"49",X"5B",X"40",X"2F",X"8F",X"2F",X"80",X"8E",X"02",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"2F",X"8F",X"2F",X"80",X"10",X"02",X"44",X"41",X"56",X"49",
		X"44",X"40",X"40",X"40",X"40",X"40",X"2F",X"81",X"2F",X"80",X"12",X"02",X"46",X"4C",X"41",X"56",
		X"49",X"41",X"40",X"40",X"40",X"40",X"2F",X"83",X"2F",X"80",X"14",X"02",X"4D",X"49",X"47",X"55",
		X"45",X"4C",X"49",X"54",X"4F",X"40",X"2F",X"85",X"2F",X"80",X"16",X"02",X"52",X"4F",X"4D",X"49",
		X"4E",X"41",X"40",X"40",X"40",X"40",X"2F",X"87",X"2F",X"80",X"18",X"02",X"4D",X"41",X"4D",X"49",
		X"40",X"40",X"40",X"40",X"40",X"40",X"2F",X"89",X"2F",X"80",X"1A",X"02",X"50",X"41",X"50",X"49",
		X"40",X"40",X"40",X"40",X"40",X"40",X"2F",X"89",X"2F",X"80",X"EF",X"00",X"01",X"EF",X"01",X"00",
		X"EF",X"04",X"00",X"EF",X"1E",X"00",X"0E",X"0C",X"CD",X"86",X"06",X"C9",X"21",X"04",X"4E",X"3E",
		X"20",X"77",X"C9",X"C9",X"F5",X"EF",X"20",X"12",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",
		X"EF",X"20",X"13",X"EF",X"21",X"12",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",X"EF",X"20",
		X"14",X"EF",X"21",X"13",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",X"EF",X"20",X"15",X"EF",
		X"21",X"14",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",X"EF",X"20",X"16",X"EF",X"21",X"15",
		X"21",X"BC",X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",X"EF",X"20",X"17",X"EF",X"21",X"16",X"21",X"BC",
		X"4E",X"CB",X"DE",X"F1",X"C9",X"F5",X"EF",X"20",X"18",X"EF",X"21",X"17",X"21",X"BC",X"4E",X"CB",
		X"DE",X"F1",X"C9",X"F5",X"EF",X"20",X"19",X"EF",X"21",X"18",X"21",X"BC",X"4E",X"CB",X"DE",X"F1",
		X"C9",X"F5",X"EF",X"20",X"1A",X"EF",X"21",X"19",X"21",X"BC",X"4E",X"CB",X"E6",X"F1",X"C9",X"3A",
		X"13",X"4E",X"3A",X"02",X"4D",X"80",X"99",X"82",X"0F",X"0F",X"0F",X"85",X"6F",X"3A",X"00",X"4D",
		X"85",X"6F",X"3A",X"04",X"4D",X"85",X"6F",X"3A",X"06",X"4D",X"85",X"E6",X"0F",X"E7",X"46",X"1D",
		X"FF",X"1C",X"22",X"1D",X"FF",X"1C",X"54",X"1D",X"1C",X"93",X"2D",X"93",X"22",X"1D",X"FF",X"1C",
		X"3E",X"93",X"22",X"1D",X"4F",X"93",X"60",X"93",X"71",X"93",X"46",X"1D",X"82",X"93",X"EF",X"7A",
		X"EF",X"7A",X"EF",X"7A",X"60",X"93",X"46",X"1D",X"FF",X"1C",X"EF",X"65",X"EF",X"7A",X"60",X"93",
		X"46",X"1D",X"FF",X"1C",X"EF",X"65",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"41",
		X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",
		X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"EF",X"A5",X"31",X"32",X"33",X"34",X"35",
		X"36",X"37",X"38",X"39",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8B",X"8C",
		X"8D",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",X"95",X"96",X"97",X"98",X"99",X"9A",X"F5",X"C5",
		X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"08",X"D9",X"F5",X"C5",X"D5",X"E5",X"21",X"00",X"60",X"11",
		X"01",X"60",X"01",X"00",X"20",X"6F",X"B7",X"ED",X"70",X"21",X"00",X"40",X"11",X"01",X"40",X"01",
		X"00",X"04",X"3E",X"80",X"ED",X"70",X"21",X"00",X"44",X"11",X"01",X"44",X"01",X"00",X"04",X"3E",
		X"0F",X"ED",X"70",X"11",X"17",X"1B",X"CD",X"6B",X"01",X"83",X"81",X"92",X"87",X"81",X"80",X"90",
		X"92",X"8F",X"87",X"92",X"81",X"8D",X"81",X"80",X"96",X"8F",X"8C",X"81",X"94",X"89",X"8C",X"00",
		X"11",X"15",X"1B",X"CD",X"6B",X"01",X"8F",X"90",X"85",X"92",X"81",X"83",X"89",X"8F",X"8E",X"80",
		X"84",X"85",X"80",X"92",X"85",X"94",X"85",X"8E",X"83",X"89",X"8F",X"8E",X"00",X"01",X"00",X"00",
		X"21",X"00",X"40",X"11",X"00",X"20",X"ED",X"B8",X"B7",X"03",X"23",X"1B",X"BB",X"72",X"20",X"F6",
		X"3E",X"0F",X"11",X"17",X"1B",X"CD",X"6B",X"01",X"90",X"92",X"8F",X"87",X"92",X"81",X"8D",X"81",
		X"80",X"96",X"8F",X"8C",X"81",X"94",X"89",X"8C",X"80",X"83",X"81",X"92",X"87",X"81",X"84",X"8F",
		X"00",X"11",X"15",X"1B",X"CD",X"6B",X"01",X"8F",X"90",X"85",X"92",X"81",X"83",X"89",X"8F",X"8E",
		X"80",X"84",X"85",X"80",X"92",X"85",X"94",X"85",X"8E",X"83",X"89",X"8F",X"8E",X"00",X"CD",X"00",
		X"60",X"CD",X"6F",X"65",X"CD",X"80",X"73",X"20",X"25",X"3E",X"0F",X"11",X"10",X"1B",X"CD",X"6B",
		X"01",X"8F",X"90",X"85",X"92",X"81",X"94",X"89",X"96",X"8F",X"80",X"8F",X"8B",X"00",X"E1",X"D1",
		X"C1",X"F1",X"D9",X"08",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"ED",X"85",X"3E",X"0F",
		X"11",X"10",X"1B",X"CD",X"6B",X"01",X"8F",X"90",X"85",X"92",X"81",X"94",X"89",X"96",X"8F",X"80",
		X"82",X"81",X"84",X"00",X"3E",X"0F",X"11",X"0E",X"1B",X"CD",X"6B",X"01",X"92",X"85",X"89",X"8E",
		X"89",X"83",X"89",X"85",X"80",X"8C",X"8F",X"81",X"84",X"80",X"8F",X"90",X"85",X"92",X"81",X"94",
		X"89",X"96",X"8F",X"00",X"E1",X"D1",X"C1",X"F1",X"D9",X"08",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",
		X"C1",X"F1",X"ED",X"85",X"1D",X"03",X"9C",X"80",X"8F",X"8A",X"85",X"84",X"81",X"80",X"31",X"39",
		X"39",X"30",X"2F",X"41",X"2F",X"40",X"85",X"03",X"80",X"26",X"80",X"80",X"84",X"8F",X"82",X"8C",
		X"85",X"80",X"80",X"83",X"8F",X"8D",X"81",X"8E",X"84",X"8F",X"80",X"80",X"27",X"80",X"2F",X"40",
		X"2F",X"40",X"85",X"03",X"80",X"26",X"80",X"80",X"84",X"8F",X"82",X"8C",X"85",X"80",X"80",X"83",
		X"8F",X"8D",X"81",X"8E",X"84",X"8F",X"80",X"80",X"27",X"80",X"2F",X"41",X"2F",X"40",X"52",X"02",
		X"80",X"80",X"94",X"95",X"92",X"82",X"8F",X"9B",X"80",X"80",X"2F",X"41",X"2F",X"40",X"52",X"02",
		X"85",X"98",X"94",X"92",X"81",X"80",X"83",X"8F",X"89",X"8E",X"2F",X"49",X"2F",X"40",X"5B",X"02",
		X"8D",X"89",X"8B",X"99",X"80",X"80",X"93",X"92",X"8C",X"2F",X"49",X"2F",X"40",X"5B",X"02",X"8D",
		X"89",X"8B",X"99",X"80",X"80",X"93",X"92",X"8C",X"2F",X"41",X"2F",X"40",X"4B",X"02",X"80",X"80",
		X"8C",X"81",X"8D",X"82",X"81",X"84",X"81",X"2F",X"45",X"2F",X"40",X"4E",X"02",X"82",X"95",X"95",
		X"95",X"95",X"9B",X"80",X"2F",X"4F",X"2F",X"40",X"10",X"02",X"8A",X"89",X"80",X"8A",X"89",X"9B",
		X"80",X"2F",X"4F",X"2F",X"40",X"4E",X"02",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"2F",X"4F",
		X"2F",X"40",X"10",X"02",X"84",X"81",X"96",X"89",X"84",X"80",X"80",X"80",X"80",X"80",X"2F",X"41",
		X"2F",X"40",X"12",X"02",X"86",X"8C",X"81",X"96",X"89",X"81",X"80",X"80",X"80",X"80",X"2F",X"43",
		X"2F",X"40",X"14",X"02",X"8D",X"89",X"87",X"95",X"85",X"8C",X"89",X"94",X"8F",X"80",X"2F",X"45",
		X"2F",X"40",X"16",X"02",X"92",X"8F",X"8D",X"89",X"8E",X"81",X"80",X"80",X"80",X"80",X"2F",X"47",
		X"2F",X"40",X"18",X"02",X"8D",X"81",X"8D",X"89",X"80",X"80",X"80",X"80",X"80",X"80",X"2F",X"49",
		X"2F",X"40",X"1A",X"02",X"90",X"81",X"90",X"89",X"80",X"80",X"80",X"80",X"80",X"80",X"2F",X"49",
		X"2F",X"40",X"CD",X"8E",X"3A",X"3E",X"0F",X"11",X"1A",X"1B",X"CD",X"6B",X"01",X"89",X"8E",X"84",
		X"95",X"93",X"94",X"92",X"89",X"81",X"80",X"81",X"92",X"87",X"85",X"8E",X"94",X"89",X"8E",X"81",
		X"00",X"06",X"10",X"CD",X"A8",X"32",X"3E",X"0F",X"11",X"1C",X"1B",X"CD",X"6B",X"01",X"9C",X"80",
		X"89",X"8E",X"87",X"80",X"8F",X"8A",X"85",X"84",X"81",X"80",X"31",X"39",X"39",X"30",X"00",X"06",
		X"10",X"CD",X"A8",X"32",X"3E",X"0F",X"11",X"1E",X"1B",X"CD",X"6B",X"01",X"8E",X"95",X"8D",X"85",
		X"92",X"8F",X"80",X"93",X"85",X"92",X"89",X"85",X"80",X"90",X"81",X"83",X"30",X"30",X"30",X"30",
		X"00",X"06",X"10",X"CD",X"A8",X"32",X"21",X"00",X"80",X"06",X"04",X"C9",X"BB",X"03",X"8E",X"8F",
		X"92",X"8D",X"81",X"8C",X"80",X"80",X"80",X"80",X"92",X"81",X"90",X"89",X"84",X"8F",X"80",X"80",
		X"80",X"80",X"94",X"95",X"92",X"82",X"8F",X"2F",X"49",X"2F",X"40",X"B8",X"03",X"80",X"80",X"80",
		X"80",X"80",X"80",X"84",X"8F",X"82",X"8C",X"85",X"80",X"83",X"8F",X"8D",X"81",X"8E",X"84",X"8F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"2F",X"49",X"2F",X"40",X"B8",X"03",X"80",X"80",X"80",X"80",
		X"80",X"80",X"84",X"8F",X"82",X"8C",X"85",X"80",X"83",X"8F",X"8D",X"81",X"8E",X"84",X"8F",X"80",
		X"80",X"80",X"80",X"80",X"80",X"2F",X"41",X"2F",X"40",X"BB",X"03",X"8E",X"8F",X"92",X"8D",X"81",
		X"8C",X"80",X"2F",X"41",X"2F",X"40",X"3B",X"02",X"92",X"81",X"90",X"89",X"84",X"8F",X"80",X"2F",
		X"41",X"2F",X"40",X"FB",X"00",X"94",X"95",X"92",X"82",X"8F",X"2F",X"41",X"2F",X"40",X"52",X"02",
		X"94",X"95",X"92",X"82",X"8F",X"2F",X"41",X"2F",X"40",X"A9",X"03",X"80",X"80",X"80",X"80",X"89",
		X"8E",X"83",X"85",X"92",X"94",X"80",X"99",X"8F",X"95",X"92",X"80",X"8E",X"81",X"8D",X"85",X"80",
		X"80",X"80",X"2F",X"49",X"2F",X"40",X"A5",X"03",X"80",X"80",X"93",X"85",X"8C",X"85",X"83",X"94",
		X"80",X"93",X"90",X"85",X"85",X"84",X"80",X"90",X"81",X"83",X"8B",X"8D",X"81",X"8E",X"2F",X"49",
		X"2F",X"40",X"BD",X"03",X"80",X"80",X"80",X"90",X"8F",X"92",X"80",X"86",X"81",X"96",X"8F",X"92",
		X"80",X"8D",X"81",X"93",X"80",X"86",X"89",X"83",X"88",X"81",X"93",X"80",X"2F",X"45",X"2F",X"40",
		X"BD",X"03",X"80",X"80",X"90",X"8F",X"92",X"80",X"86",X"81",X"96",X"8F",X"92",X"80",X"93",X"85",
		X"8C",X"85",X"83",X"83",X"89",X"8F",X"8E",X"85",X"80",X"80",X"2F",X"45",X"2F",X"40",X"52",X"02",
		X"85",X"98",X"94",X"92",X"81",X"80",X"8C",X"89",X"86",X"85",X"2F",X"49",X"2F",X"40",X"52",X"02",
		X"82",X"8F",X"8E",X"95",X"93",X"80",X"8E",X"8F",X"8E",X"85",X"2F",X"41",X"2F",X"40",X"52",X"02",
		X"32",X"30",X"30",X"80",X"80",X"82",X"8F",X"8E",X"95",X"93",X"2F",X"45",X"2F",X"40",X"52",X"02",
		X"33",X"30",X"30",X"80",X"80",X"82",X"8F",X"8E",X"95",X"93",X"2F",X"45",X"2F",X"40",X"52",X"02",
		X"34",X"30",X"30",X"80",X"80",X"82",X"8F",X"8E",X"95",X"93",X"2F",X"45",X"2F",X"40",X"52",X"02",
		X"35",X"30",X"30",X"80",X"80",X"82",X"8F",X"8E",X"95",X"93",X"2F",X"45",X"2F",X"40",X"52",X"02",
		X"36",X"30",X"30",X"80",X"80",X"82",X"8F",X"8E",X"95",X"93",X"2F",X"45",X"2F",X"40",X"52",X"02",
		X"37",X"30",X"30",X"80",X"80",X"82",X"8F",X"8E",X"95",X"93",X"2F",X"45",X"2F",X"40",X"52",X"02",
		X"38",X"30",X"30",X"80",X"80",X"82",X"8F",X"8E",X"95",X"93",X"2F",X"45",X"2F",X"40",X"52",X"02",
		X"35",X"30",X"30",X"30",X"80",X"82",X"8F",X"8E",X"95",X"93",X"2F",X"45",X"2F",X"40",X"D4",X"43",
		X"8D",X"89",X"8B",X"99",X"80",X"83",X"88",X"85",X"8C",X"8F",X"2F",X"41",X"2F",X"40",X"4C",X"02",
		X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"2F",X"45",X"2F",X"40",X"3B",X"40",
		X"83",X"92",X"85",X"84",X"89",X"94",X"80",X"80",X"80",X"2F",X"4F",X"2F",X"40",X"3B",X"40",X"86",
		X"92",X"85",X"85",X"80",X"90",X"8C",X"81",X"99",X"2F",X"4F",X"2F",X"40",X"4C",X"02",X"90",X"8C",
		X"81",X"99",X"85",X"92",X"80",X"8F",X"8E",X"85",X"2F",X"45",X"4C",X"02",X"90",X"8C",X"81",X"99",
		X"85",X"92",X"80",X"94",X"97",X"8F",X"2F",X"45",X"2F",X"40",X"52",X"02",X"87",X"81",X"8D",X"85",
		X"80",X"80",X"8F",X"96",X"85",X"92",X"2F",X"41",X"2F",X"40",X"92",X"02",X"92",X"85",X"81",X"84",
		X"99",X"9B",X"2F",X"49",X"2F",X"50",X"ED",X"02",X"90",X"95",X"93",X"88",X"80",X"93",X"94",X"81",
		X"92",X"94",X"80",X"82",X"95",X"94",X"94",X"8F",X"8E",X"2F",X"47",X"2F",X"40",X"6F",X"02",X"31",
		X"80",X"90",X"8C",X"81",X"99",X"85",X"92",X"80",X"8F",X"8E",X"8C",X"99",X"80",X"2F",X"47",X"2F",
		X"40",X"6F",X"02",X"31",X"80",X"8F",X"92",X"80",X"32",X"80",X"90",X"8C",X"81",X"99",X"85",X"92",
		X"93",X"2F",X"47",X"00",X"2F",X"00",X"40",X"00",X"71",X"02",X"32",X"80",X"8F",X"92",X"80",X"34",
		X"80",X"90",X"8C",X"81",X"99",X"85",X"92",X"93",X"2F",X"47",X"00",X"2F",X"00",X"40",X"00",X"56",
		X"03",X"82",X"8F",X"8E",X"95",X"93",X"80",X"90",X"95",X"83",X"8B",X"8D",X"81",X"8E",X"80",X"86",
		X"8F",X"92",X"80",X"80",X"80",X"30",X"30",X"30",X"80",X"9D",X"9E",X"9F",X"2F",X"4E",X"2F",X"40",
		X"04",X"03",X"8D",X"85",X"8D",X"8F",X"92",X"99",X"80",X"80",X"8F",X"8B",X"2F",X"4F",X"2F",X"40",
		X"04",X"03",X"82",X"81",X"84",X"80",X"80",X"80",X"80",X"92",X"80",X"8D",X"2F",X"4F",X"2F",X"40",
		X"08",X"03",X"31",X"80",X"83",X"8F",X"89",X"8E",X"80",X"80",X"31",X"80",X"83",X"92",X"85",X"84",
		X"89",X"94",X"80",X"2F",X"4F",X"2F",X"40",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"95",
		X"95",X"95",X"95",X"95",X"95",X"84",X"85",X"93",X"81",X"92",X"92",X"8F",X"8C",X"8C",X"8F",X"20",
		X"84",X"85",X"8C",X"20",X"89",X"8E",X"87",X"85",X"8E",X"89",X"85",X"92",X"8F",X"20",X"8D",X"89",
		X"87",X"95",X"85",X"8C",X"20",X"81",X"8E",X"94",X"8F",X"8E",X"89",X"8F",X"20",X"8F",X"8A",X"85",
		X"84",X"81",X"20",X"20",X"92",X"85",X"81",X"8C",X"89",X"9A",X"81",X"84",X"8F",X"20",X"85",X"8C",
		X"20",X"31",X"30",X"2F",X"31",X"32",X"2F",X"38",X"39",X"20",X"93",X"8F",X"82",X"92",X"85",X"20",
		X"95",X"8E",X"81",X"20",X"90",X"8C",X"81",X"83",X"81",X"20",X"84",X"85",X"20",X"8D",X"93",X"93",
		X"20",X"20",X"20",X"90",X"81",X"83",X"8B",X"8D",X"81",X"8E",X"20",X"90",X"81",X"92",X"81",X"20",
		X"8D",X"85",X"8A",X"8F",X"92",X"81",X"92",X"20",X"8C",X"81",X"20",X"90",X"85",X"92",X"86",X"8F",
		X"8D",X"81",X"8E",X"93",X"20",X"84",X"85",X"20",X"85",X"93",X"94",X"81",X"20",X"20",X"20",X"20",
		X"20",X"20",X"81",X"94",X"85",X"8E",X"83",X"89",X"8F",X"8E",X"3A",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"85",X"8E",X"20",X"83",X"81",X"93",X"8F",X"20",X"84",X"85",X"20",
		X"94",X"85",X"8E",X"85",X"92",X"20",X"95",X"8E",X"81",X"20",X"90",X"85",X"92",X"84",X"89",X"84",
		X"81",X"20",X"84",X"85",X"8C",X"20",X"93",X"89",X"93",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"90",X"8F",X"8E",X"85",X"92",X"93",X"85",X"20",X"85",X"8E",X"20",X"83",X"8F",X"8E",X"94",X"81",
		X"83",X"94",X"8F",X"20",X"83",X"8F",X"8E",X"20",X"8D",X"89",X"8B",X"99",X"20",X"93",X"2E",X"92",
		X"2E",X"8C",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"83",
		X"8F",X"84",X"89",X"87",X"8F",X"20",X"90",X"8F",X"93",X"94",X"81",X"8C",X"20",X"31",X"34",X"30",
		X"37",X"20",X"81",X"92",X"81",X"8E",X"87",X"95",X"92",X"85",X"8E",X"20",X"34",X"31",X"34",X"38",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"83",X"81",
		X"90",X"89",X"94",X"81",X"8C",X"20",X"86",X"85",X"84",X"85",X"92",X"81",X"8C",X"20",X"92",X"85",
		X"90",X"95",X"82",X"8C",X"89",X"83",X"81",X"20",X"81",X"92",X"87",X"85",X"8E",X"94",X"89",X"8E",
		X"81",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"94",X"85",X"8C",
		X"20",X"36",X"39",X"2D",X"39",X"38",X"35",X"31",X"20",X"36",X"37",X"2D",X"39",X"33",X"38",X"33",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"95",X"8E",X"81",X"20",X"8D",X"81",X"8E",X"89",X"90",X"95",X"8C",X"81",X"83",X"89",X"8F",X"8E",
		X"20",X"89",X"8E",X"84",X"85",X"96",X"89",X"84",X"81",X"20",X"83",X"81",X"8E",X"83",X"85",X"8C",
		X"81",X"20",X"8C",X"81",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"87",X"81",X"92",X"81",X"8E",
		X"94",X"89",X"81",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"88",X"85",X"83",X"88",X"8F",X"20",X"85",
		X"8C",X"20",X"84",X"85",X"90",X"8F",X"93",X"89",X"94",X"8F",X"20",X"91",X"95",X"85",X"20",X"8D",
		X"81",X"92",X"83",X"81",X"20",X"8C",X"81",X"20",X"8C",X"85",X"99",X"20",X"31",X"31",X"37",X"32",
		X"33",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"91",X"95",X"85",X"84",X"81",X"20",X"92",X"85",
		X"87",X"89",X"93",X"94",X"92",X"81",X"84",X"8F",X"20",X"85",X"8E",X"20",X"94",X"85",X"92",X"92",
		X"89",X"94",X"8F",X"92",X"89",X"8F",X"20",X"84",X"85",X"20",X"8C",X"81",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"92",X"85",X"90",X"95",X"82",X"8C",X"89",X"83",X"81",
		X"20",X"81",X"92",X"87",X"85",X"8E",X"94",X"89",X"8E",X"81",X"20",X"85",X"8C",X"20",X"93",X"8F",
		X"86",X"94",X"97",X"81",X"92",X"85",X"20",X"83",X"8C",X"95",X"82",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"83",X"95",X"81",X"8C",X"91",X"95",X"89",X"85",X"92",X"20",
		X"92",X"85",X"90",X"92",X"8F",X"84",X"95",X"83",X"83",X"89",X"8F",X"8E",X"20",X"90",X"81",X"92",
		X"83",X"89",X"81",X"8C",X"20",X"99",X"2F",X"8F",X"20",X"94",X"8F",X"94",X"81",X"8C",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"84",X"85",X"20",X"85",X"93",X"94",X"81",X"20",X"93",X"85",X"92",
		X"81",X"20",X"90",X"85",X"8E",X"81",X"84",X"81",X"20",X"83",X"8F",X"8E",X"20",X"8C",X"8F",X"93",
		X"20",X"81",X"8C",X"83",X"81",X"8E",X"83",X"85",X"93",X"20",X"84",X"85",X"20",X"8C",X"81",X"20",
		X"20",X"20",X"20",X"20",X"8C",X"85",X"99",X"20",X"31",X"31",X"37",X"32",X"33",X"20",X"2E",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"E5",
		X"F5",X"2A",X"6C",X"4C",X"7D",X"B4",X"28",X"03",X"F1",X"E1",X"C9",X"F1",X"3E",X"F3",X"E1",X"C9");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
